library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LED_Flash_LUT_pkg is
 
 type my_array is array (4095 downto 0) of integer;
 constant DtoP_LUT : my_array := (
 
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	60000	)	,
(	59983	)	,
(	59966	)	,
(	59949	)	,
(	59932	)	,
(	59915	)	,
(	59898	)	,
(	59881	)	,
(	59864	)	,
(	59847	)	,
(	59830	)	,
(	59813	)	,
(	59796	)	,
(	59779	)	,
(	59762	)	,
(	59745	)	,
(	59728	)	,
(	59711	)	,
(	59694	)	,
(	59677	)	,
(	59660	)	,
(	59643	)	,
(	59626	)	,
(	59609	)	,
(	59592	)	,
(	59575	)	,
(	59558	)	,
(	59541	)	,
(	59524	)	,
(	59507	)	,
(	59490	)	,
(	59473	)	,
(	59456	)	,
(	59439	)	,
(	59422	)	,
(	59405	)	,
(	59388	)	,
(	59371	)	,
(	59354	)	,
(	59337	)	,
(	59320	)	,
(	59303	)	,
(	59286	)	,
(	59269	)	,
(	59252	)	,
(	59235	)	,
(	59218	)	,
(	59201	)	,
(	59184	)	,
(	59167	)	,
(	59150	)	,
(	59133	)	,
(	59116	)	,
(	59099	)	,
(	59082	)	,
(	59065	)	,
(	59048	)	,
(	59031	)	,
(	59014	)	,
(	58997	)	,
(	58980	)	,
(	58963	)	,
(	58946	)	,
(	58929	)	,
(	58912	)	,
(	58895	)	,
(	58878	)	,
(	58861	)	,
(	58844	)	,
(	58827	)	,
(	58810	)	,
(	58793	)	,
(	58776	)	,
(	58759	)	,
(	58742	)	,
(	58725	)	,
(	58708	)	,
(	58691	)	,
(	58674	)	,
(	58657	)	,
(	58640	)	,
(	58623	)	,
(	58606	)	,
(	58589	)	,
(	58572	)	,
(	58555	)	,
(	58538	)	,
(	58521	)	,
(	58504	)	,
(	58487	)	,
(	58470	)	,
(	58453	)	,
(	58436	)	,
(	58419	)	,
(	58402	)	,
(	58385	)	,
(	58368	)	,
(	58351	)	,
(	58334	)	,
(	58317	)	,
(	58300	)	,
(	58283	)	,
(	58266	)	,
(	58249	)	,
(	58232	)	,
(	58215	)	,
(	58198	)	,
(	58181	)	,
(	58164	)	,
(	58147	)	,
(	58130	)	,
(	58113	)	,
(	58096	)	,
(	58079	)	,
(	58062	)	,
(	58045	)	,
(	58028	)	,
(	58011	)	,
(	57994	)	,
(	57977	)	,
(	57960	)	,
(	57943	)	,
(	57926	)	,
(	57909	)	,
(	57892	)	,
(	57875	)	,
(	57858	)	,
(	57841	)	,
(	57824	)	,
(	57807	)	,
(	57790	)	,
(	57773	)	,
(	57756	)	,
(	57739	)	,
(	57722	)	,
(	57705	)	,
(	57688	)	,
(	57671	)	,
(	57654	)	,
(	57637	)	,
(	57620	)	,
(	57603	)	,
(	57586	)	,
(	57569	)	,
(	57552	)	,
(	57535	)	,
(	57518	)	,
(	57501	)	,
(	57484	)	,
(	57467	)	,
(	57450	)	,
(	57433	)	,
(	57416	)	,
(	57399	)	,
(	57382	)	,
(	57365	)	,
(	57348	)	,
(	57331	)	,
(	57314	)	,
(	57297	)	,
(	57280	)	,
(	57263	)	,
(	57246	)	,
(	57229	)	,
(	57212	)	,
(	57195	)	,
(	57178	)	,
(	57161	)	,
(	57144	)	,
(	57127	)	,
(	57110	)	,
(	57093	)	,
(	57076	)	,
(	57059	)	,
(	57042	)	,
(	57025	)	,
(	57008	)	,
(	56991	)	,
(	56974	)	,
(	56957	)	,
(	56940	)	,
(	56923	)	,
(	56906	)	,
(	56889	)	,
(	56872	)	,
(	56855	)	,
(	56838	)	,
(	56821	)	,
(	56804	)	,
(	56787	)	,
(	56770	)	,
(	56753	)	,
(	56736	)	,
(	56719	)	,
(	56702	)	,
(	56685	)	,
(	56668	)	,
(	56651	)	,
(	56634	)	,
(	56617	)	,
(	56600	)	,
(	56583	)	,
(	56566	)	,
(	56549	)	,
(	56532	)	,
(	56515	)	,
(	56498	)	,
(	56481	)	,
(	56464	)	,
(	56447	)	,
(	56430	)	,
(	56413	)	,
(	56396	)	,
(	56379	)	,
(	56362	)	,
(	56345	)	,
(	56328	)	,
(	56311	)	,
(	56294	)	,
(	56277	)	,
(	56260	)	,
(	56243	)	,
(	56226	)	,
(	56209	)	,
(	56192	)	,
(	56175	)	,
(	56158	)	,
(	56141	)	,
(	56124	)	,
(	56107	)	,
(	56090	)	,
(	56073	)	,
(	56056	)	,
(	56039	)	,
(	56022	)	,
(	56005	)	,
(	55988	)	,
(	55971	)	,
(	55954	)	,
(	55937	)	,
(	55920	)	,
(	55903	)	,
(	55886	)	,
(	55869	)	,
(	55852	)	,
(	55835	)	,
(	55818	)	,
(	55801	)	,
(	55784	)	,
(	55767	)	,
(	55750	)	,
(	55733	)	,
(	55716	)	,
(	55699	)	,
(	55682	)	,
(	55665	)	,
(	55648	)	,
(	55631	)	,
(	55614	)	,
(	55597	)	,
(	55580	)	,
(	55563	)	,
(	55546	)	,
(	55529	)	,
(	55512	)	,
(	55495	)	,
(	55478	)	,
(	55461	)	,
(	55444	)	,
(	55427	)	,
(	55410	)	,
(	55393	)	,
(	55376	)	,
(	55359	)	,
(	55342	)	,
(	55325	)	,
(	55308	)	,
(	55291	)	,
(	55274	)	,
(	55257	)	,
(	55240	)	,
(	55223	)	,
(	55206	)	,
(	55189	)	,
(	55172	)	,
(	55155	)	,
(	55138	)	,
(	55121	)	,
(	55104	)	,
(	55087	)	,
(	55070	)	,
(	55053	)	,
(	55036	)	,
(	55019	)	,
(	55002	)	,
(	54985	)	,
(	54968	)	,
(	54951	)	,
(	54934	)	,
(	54917	)	,
(	54900	)	,
(	54883	)	,
(	54866	)	,
(	54849	)	,
(	54832	)	,
(	54815	)	,
(	54798	)	,
(	54781	)	,
(	54764	)	,
(	54747	)	,
(	54730	)	,
(	54713	)	,
(	54696	)	,
(	54679	)	,
(	54662	)	,
(	54645	)	,
(	54628	)	,
(	54611	)	,
(	54594	)	,
(	54577	)	,
(	54560	)	,
(	54543	)	,
(	54526	)	,
(	54509	)	,
(	54492	)	,
(	54475	)	,
(	54458	)	,
(	54441	)	,
(	54424	)	,
(	54407	)	,
(	54390	)	,
(	54373	)	,
(	54356	)	,
(	54339	)	,
(	54322	)	,
(	54305	)	,
(	54288	)	,
(	54271	)	,
(	54254	)	,
(	54237	)	,
(	54220	)	,
(	54203	)	,
(	54186	)	,
(	54169	)	,
(	54152	)	,
(	54135	)	,
(	54118	)	,
(	54101	)	,
(	54084	)	,
(	54067	)	,
(	54050	)	,
(	54033	)	,
(	54016	)	,
(	53999	)	,
(	53982	)	,
(	53965	)	,
(	53948	)	,
(	53931	)	,
(	53914	)	,
(	53897	)	,
(	53880	)	,
(	53863	)	,
(	53846	)	,
(	53829	)	,
(	53812	)	,
(	53795	)	,
(	53778	)	,
(	53761	)	,
(	53744	)	,
(	53727	)	,
(	53710	)	,
(	53693	)	,
(	53676	)	,
(	53659	)	,
(	53642	)	,
(	53625	)	,
(	53608	)	,
(	53591	)	,
(	53574	)	,
(	53557	)	,
(	53540	)	,
(	53523	)	,
(	53506	)	,
(	53489	)	,
(	53472	)	,
(	53455	)	,
(	53438	)	,
(	53421	)	,
(	53404	)	,
(	53387	)	,
(	53370	)	,
(	53353	)	,
(	53336	)	,
(	53319	)	,
(	53302	)	,
(	53285	)	,
(	53268	)	,
(	53251	)	,
(	53234	)	,
(	53217	)	,
(	53200	)	,
(	53183	)	,
(	53166	)	,
(	53149	)	,
(	53132	)	,
(	53115	)	,
(	53098	)	,
(	53081	)	,
(	53064	)	,
(	53047	)	,
(	53030	)	,
(	53013	)	,
(	52996	)	,
(	52979	)	,
(	52962	)	,
(	52945	)	,
(	52928	)	,
(	52911	)	,
(	52894	)	,
(	52877	)	,
(	52860	)	,
(	52843	)	,
(	52826	)	,
(	52809	)	,
(	52792	)	,
(	52775	)	,
(	52758	)	,
(	52741	)	,
(	52724	)	,
(	52707	)	,
(	52690	)	,
(	52673	)	,
(	52656	)	,
(	52639	)	,
(	52622	)	,
(	52605	)	,
(	52588	)	,
(	52571	)	,
(	52554	)	,
(	52537	)	,
(	52520	)	,
(	52503	)	,
(	52486	)	,
(	52469	)	,
(	52452	)	,
(	52435	)	,
(	52418	)	,
(	52401	)	,
(	52384	)	,
(	52367	)	,
(	52350	)	,
(	52333	)	,
(	52316	)	,
(	52299	)	,
(	52282	)	,
(	52265	)	,
(	52248	)	,
(	52231	)	,
(	52214	)	,
(	52197	)	,
(	52180	)	,
(	52163	)	,
(	52146	)	,
(	52129	)	,
(	52112	)	,
(	52095	)	,
(	52078	)	,
(	52061	)	,
(	52044	)	,
(	52027	)	,
(	52010	)	,
(	51993	)	,
(	51976	)	,
(	51959	)	,
(	51942	)	,
(	51925	)	,
(	51908	)	,
(	51891	)	,
(	51874	)	,
(	51857	)	,
(	51840	)	,
(	51823	)	,
(	51806	)	,
(	51789	)	,
(	51772	)	,
(	51755	)	,
(	51738	)	,
(	51721	)	,
(	51704	)	,
(	51687	)	,
(	51670	)	,
(	51653	)	,
(	51636	)	,
(	51619	)	,
(	51602	)	,
(	51585	)	,
(	51568	)	,
(	51551	)	,
(	51534	)	,
(	51517	)	,
(	51500	)	,
(	51483	)	,
(	51466	)	,
(	51449	)	,
(	51432	)	,
(	51415	)	,
(	51398	)	,
(	51381	)	,
(	51364	)	,
(	51347	)	,
(	51330	)	,
(	51313	)	,
(	51296	)	,
(	51279	)	,
(	51262	)	,
(	51245	)	,
(	51228	)	,
(	51211	)	,
(	51194	)	,
(	51177	)	,
(	51160	)	,
(	51143	)	,
(	51126	)	,
(	51109	)	,
(	51092	)	,
(	51075	)	,
(	51058	)	,
(	51041	)	,
(	51024	)	,
(	51007	)	,
(	50990	)	,
(	50973	)	,
(	50956	)	,
(	50939	)	,
(	50922	)	,
(	50905	)	,
(	50888	)	,
(	50871	)	,
(	50854	)	,
(	50837	)	,
(	50820	)	,
(	50803	)	,
(	50786	)	,
(	50769	)	,
(	50752	)	,
(	50735	)	,
(	50718	)	,
(	50701	)	,
(	50684	)	,
(	50667	)	,
(	50650	)	,
(	50633	)	,
(	50616	)	,
(	50599	)	,
(	50582	)	,
(	50565	)	,
(	50548	)	,
(	50531	)	,
(	50514	)	,
(	50497	)	,
(	50480	)	,
(	50463	)	,
(	50446	)	,
(	50429	)	,
(	50412	)	,
(	50395	)	,
(	50378	)	,
(	50361	)	,
(	50344	)	,
(	50327	)	,
(	50310	)	,
(	50293	)	,
(	50276	)	,
(	50259	)	,
(	50242	)	,
(	50225	)	,
(	50208	)	,
(	50191	)	,
(	50174	)	,
(	50157	)	,
(	50140	)	,
(	50123	)	,
(	50106	)	,
(	50089	)	,
(	50072	)	,
(	50055	)	,
(	50038	)	,
(	50021	)	,
(	50004	)	,
(	49987	)	,
(	49970	)	,
(	49953	)	,
(	49936	)	,
(	49919	)	,
(	49902	)	,
(	49885	)	,
(	49868	)	,
(	49851	)	,
(	49834	)	,
(	49817	)	,
(	49800	)	,
(	49783	)	,
(	49766	)	,
(	49749	)	,
(	49732	)	,
(	49715	)	,
(	49698	)	,
(	49681	)	,
(	49664	)	,
(	49647	)	,
(	49630	)	,
(	49613	)	,
(	49596	)	,
(	49579	)	,
(	49562	)	,
(	49545	)	,
(	49528	)	,
(	49511	)	,
(	49494	)	,
(	49477	)	,
(	49460	)	,
(	49443	)	,
(	49426	)	,
(	49409	)	,
(	49392	)	,
(	49375	)	,
(	49358	)	,
(	49341	)	,
(	49324	)	,
(	49307	)	,
(	49290	)	,
(	49273	)	,
(	49256	)	,
(	49239	)	,
(	49222	)	,
(	49205	)	,
(	49188	)	,
(	49171	)	,
(	49154	)	,
(	49137	)	,
(	49120	)	,
(	49103	)	,
(	49086	)	,
(	49069	)	,
(	49052	)	,
(	49035	)	,
(	49018	)	,
(	49001	)	,
(	48984	)	,
(	48967	)	,
(	48950	)	,
(	48933	)	,
(	48916	)	,
(	48899	)	,
(	48882	)	,
(	48865	)	,
(	48848	)	,
(	48831	)	,
(	48814	)	,
(	48797	)	,
(	48780	)	,
(	48763	)	,
(	48746	)	,
(	48729	)	,
(	48712	)	,
(	48695	)	,
(	48678	)	,
(	48661	)	,
(	48644	)	,
(	48627	)	,
(	48610	)	,
(	48593	)	,
(	48576	)	,
(	48559	)	,
(	48542	)	,
(	48525	)	,
(	48508	)	,
(	48491	)	,
(	48474	)	,
(	48457	)	,
(	48440	)	,
(	48423	)	,
(	48406	)	,
(	48389	)	,
(	48372	)	,
(	48355	)	,
(	48338	)	,
(	48321	)	,
(	48304	)	,
(	48287	)	,
(	48270	)	,
(	48253	)	,
(	48236	)	,
(	48219	)	,
(	48202	)	,
(	48185	)	,
(	48168	)	,
(	48151	)	,
(	48134	)	,
(	48117	)	,
(	48100	)	,
(	48083	)	,
(	48066	)	,
(	48049	)	,
(	48032	)	,
(	48015	)	,
(	47998	)	,
(	47981	)	,
(	47964	)	,
(	47947	)	,
(	47930	)	,
(	47913	)	,
(	47896	)	,
(	47879	)	,
(	47862	)	,
(	47845	)	,
(	47828	)	,
(	47811	)	,
(	47794	)	,
(	47777	)	,
(	47760	)	,
(	47743	)	,
(	47726	)	,
(	47709	)	,
(	47692	)	,
(	47675	)	,
(	47658	)	,
(	47641	)	,
(	47624	)	,
(	47607	)	,
(	47590	)	,
(	47573	)	,
(	47556	)	,
(	47539	)	,
(	47522	)	,
(	47505	)	,
(	47488	)	,
(	47471	)	,
(	47454	)	,
(	47437	)	,
(	47420	)	,
(	47403	)	,
(	47386	)	,
(	47369	)	,
(	47352	)	,
(	47335	)	,
(	47318	)	,
(	47301	)	,
(	47284	)	,
(	47267	)	,
(	47250	)	,
(	47233	)	,
(	47216	)	,
(	47199	)	,
(	47182	)	,
(	47165	)	,
(	47148	)	,
(	47131	)	,
(	47114	)	,
(	47097	)	,
(	47080	)	,
(	47063	)	,
(	47046	)	,
(	47029	)	,
(	47012	)	,
(	46995	)	,
(	46978	)	,
(	46961	)	,
(	46944	)	,
(	46927	)	,
(	46910	)	,
(	46893	)	,
(	46876	)	,
(	46859	)	,
(	46842	)	,
(	46825	)	,
(	46808	)	,
(	46791	)	,
(	46774	)	,
(	46757	)	,
(	46740	)	,
(	46723	)	,
(	46706	)	,
(	46689	)	,
(	46672	)	,
(	46655	)	,
(	46638	)	,
(	46621	)	,
(	46604	)	,
(	46587	)	,
(	46570	)	,
(	46553	)	,
(	46536	)	,
(	46519	)	,
(	46502	)	,
(	46485	)	,
(	46468	)	,
(	46451	)	,
(	46434	)	,
(	46417	)	,
(	46400	)	,
(	46383	)	,
(	46366	)	,
(	46349	)	,
(	46332	)	,
(	46315	)	,
(	46298	)	,
(	46281	)	,
(	46264	)	,
(	46247	)	,
(	46230	)	,
(	46213	)	,
(	46196	)	,
(	46179	)	,
(	46162	)	,
(	46145	)	,
(	46128	)	,
(	46111	)	,
(	46094	)	,
(	46077	)	,
(	46060	)	,
(	46043	)	,
(	46026	)	,
(	46009	)	,
(	45992	)	,
(	45975	)	,
(	45958	)	,
(	45941	)	,
(	45924	)	,
(	45907	)	,
(	45890	)	,
(	45873	)	,
(	45856	)	,
(	45839	)	,
(	45822	)	,
(	45805	)	,
(	45788	)	,
(	45771	)	,
(	45754	)	,
(	45737	)	,
(	45720	)	,
(	45703	)	,
(	45686	)	,
(	45669	)	,
(	45652	)	,
(	45635	)	,
(	45618	)	,
(	45601	)	,
(	45584	)	,
(	45567	)	,
(	45550	)	,
(	45533	)	,
(	45516	)	,
(	45499	)	,
(	45482	)	,
(	45465	)	,
(	45448	)	,
(	45431	)	,
(	45414	)	,
(	45397	)	,
(	45380	)	,
(	45363	)	,
(	45346	)	,
(	45329	)	,
(	45312	)	,
(	45295	)	,
(	45278	)	,
(	45261	)	,
(	45244	)	,
(	45227	)	,
(	45210	)	,
(	45193	)	,
(	45176	)	,
(	45159	)	,
(	45142	)	,
(	45125	)	,
(	45108	)	,
(	45091	)	,
(	45074	)	,
(	45057	)	,
(	45040	)	,
(	45023	)	,
(	45006	)	,
(	44989	)	,
(	44972	)	,
(	44955	)	,
(	44938	)	,
(	44921	)	,
(	44904	)	,
(	44887	)	,
(	44870	)	,
(	44853	)	,
(	44836	)	,
(	44819	)	,
(	44802	)	,
(	44785	)	,
(	44768	)	,
(	44751	)	,
(	44734	)	,
(	44717	)	,
(	44700	)	,
(	44683	)	,
(	44666	)	,
(	44649	)	,
(	44632	)	,
(	44615	)	,
(	44598	)	,
(	44581	)	,
(	44564	)	,
(	44547	)	,
(	44530	)	,
(	44513	)	,
(	44496	)	,
(	44479	)	,
(	44462	)	,
(	44445	)	,
(	44428	)	,
(	44411	)	,
(	44394	)	,
(	44377	)	,
(	44360	)	,
(	44343	)	,
(	44326	)	,
(	44309	)	,
(	44292	)	,
(	44275	)	,
(	44258	)	,
(	44241	)	,
(	44224	)	,
(	44207	)	,
(	44190	)	,
(	44173	)	,
(	44156	)	,
(	44139	)	,
(	44122	)	,
(	44105	)	,
(	44088	)	,
(	44071	)	,
(	44054	)	,
(	44037	)	,
(	44020	)	,
(	44003	)	,
(	43986	)	,
(	43969	)	,
(	43952	)	,
(	43935	)	,
(	43918	)	,
(	43901	)	,
(	43884	)	,
(	43867	)	,
(	43850	)	,
(	43833	)	,
(	43816	)	,
(	43799	)	,
(	43782	)	,
(	43765	)	,
(	43748	)	,
(	43731	)	,
(	43714	)	,
(	43697	)	,
(	43680	)	,
(	43663	)	,
(	43646	)	,
(	43629	)	,
(	43612	)	,
(	43595	)	,
(	43578	)	,
(	43561	)	,
(	43544	)	,
(	43527	)	,
(	43510	)	,
(	43493	)	,
(	43476	)	,
(	43459	)	,
(	43442	)	,
(	43425	)	,
(	43408	)	,
(	43391	)	,
(	43374	)	,
(	43357	)	,
(	43340	)	,
(	43323	)	,
(	43306	)	,
(	43289	)	,
(	43272	)	,
(	43255	)	,
(	43238	)	,
(	43221	)	,
(	43204	)	,
(	43187	)	,
(	43170	)	,
(	43153	)	,
(	43136	)	,
(	43119	)	,
(	43102	)	,
(	43085	)	,
(	43068	)	,
(	43051	)	,
(	43034	)	,
(	43017	)	,
(	43000	)	,
(	42983	)	,
(	42966	)	,
(	42949	)	,
(	42932	)	,
(	42915	)	,
(	42898	)	,
(	42881	)	,
(	42864	)	,
(	42847	)	,
(	42830	)	,
(	42813	)	,
(	42796	)	,
(	42779	)	,
(	42762	)	,
(	42745	)	,
(	42728	)	,
(	42711	)	,
(	42694	)	,
(	42677	)	,
(	42660	)	,
(	42643	)	,
(	42626	)	,
(	42609	)	,
(	42592	)	,
(	42575	)	,
(	42558	)	,
(	42541	)	,
(	42524	)	,
(	42507	)	,
(	42490	)	,
(	42473	)	,
(	42456	)	,
(	42439	)	,
(	42422	)	,
(	42405	)	,
(	42388	)	,
(	42371	)	,
(	42354	)	,
(	42337	)	,
(	42320	)	,
(	42303	)	,
(	42286	)	,
(	42269	)	,
(	42252	)	,
(	42235	)	,
(	42218	)	,
(	42201	)	,
(	42184	)	,
(	42167	)	,
(	42150	)	,
(	42133	)	,
(	42116	)	,
(	42099	)	,
(	42082	)	,
(	42065	)	,
(	42048	)	,
(	42031	)	,
(	42014	)	,
(	41997	)	,
(	41980	)	,
(	41963	)	,
(	41946	)	,
(	41929	)	,
(	41912	)	,
(	41895	)	,
(	41878	)	,
(	41861	)	,
(	41844	)	,
(	41827	)	,
(	41810	)	,
(	41793	)	,
(	41776	)	,
(	41759	)	,
(	41742	)	,
(	41725	)	,
(	41708	)	,
(	41691	)	,
(	41674	)	,
(	41657	)	,
(	41640	)	,
(	41623	)	,
(	41606	)	,
(	41589	)	,
(	41572	)	,
(	41555	)	,
(	41538	)	,
(	41521	)	,
(	41504	)	,
(	41487	)	,
(	41470	)	,
(	41453	)	,
(	41436	)	,
(	41419	)	,
(	41402	)	,
(	41385	)	,
(	41368	)	,
(	41351	)	,
(	41334	)	,
(	41317	)	,
(	41300	)	,
(	41283	)	,
(	41266	)	,
(	41249	)	,
(	41232	)	,
(	41215	)	,
(	41198	)	,
(	41181	)	,
(	41164	)	,
(	41147	)	,
(	41130	)	,
(	41113	)	,
(	41096	)	,
(	41079	)	,
(	41062	)	,
(	41045	)	,
(	41028	)	,
(	41011	)	,
(	40994	)	,
(	40977	)	,
(	40960	)	,
(	40943	)	,
(	40926	)	,
(	40909	)	,
(	40892	)	,
(	40875	)	,
(	40858	)	,
(	40841	)	,
(	40824	)	,
(	40807	)	,
(	40790	)	,
(	40773	)	,
(	40756	)	,
(	40739	)	,
(	40722	)	,
(	40705	)	,
(	40688	)	,
(	40671	)	,
(	40654	)	,
(	40637	)	,
(	40620	)	,
(	40603	)	,
(	40586	)	,
(	40569	)	,
(	40552	)	,
(	40535	)	,
(	40518	)	,
(	40501	)	,
(	40484	)	,
(	40467	)	,
(	40450	)	,
(	40433	)	,
(	40416	)	,
(	40399	)	,
(	40382	)	,
(	40365	)	,
(	40348	)	,
(	40331	)	,
(	40314	)	,
(	40297	)	,
(	40280	)	,
(	40263	)	,
(	40246	)	,
(	40229	)	,
(	40212	)	,
(	40195	)	,
(	40178	)	,
(	40161	)	,
(	40144	)	,
(	40127	)	,
(	40110	)	,
(	40093	)	,
(	40076	)	,
(	40059	)	,
(	40042	)	,
(	40025	)	,
(	40008	)	,
(	39991	)	,
(	39974	)	,
(	39957	)	,
(	39940	)	,
(	39923	)	,
(	39906	)	,
(	39889	)	,
(	39872	)	,
(	39855	)	,
(	39838	)	,
(	39821	)	,
(	39804	)	,
(	39787	)	,
(	39770	)	,
(	39753	)	,
(	39736	)	,
(	39719	)	,
(	39702	)	,
(	39685	)	,
(	39668	)	,
(	39651	)	,
(	39634	)	,
(	39617	)	,
(	39600	)	,
(	39583	)	,
(	39566	)	,
(	39549	)	,
(	39532	)	,
(	39515	)	,
(	39498	)	,
(	39481	)	,
(	39464	)	,
(	39447	)	,
(	39430	)	,
(	39413	)	,
(	39396	)	,
(	39379	)	,
(	39362	)	,
(	39345	)	,
(	39328	)	,
(	39311	)	,
(	39294	)	,
(	39277	)	,
(	39260	)	,
(	39243	)	,
(	39226	)	,
(	39209	)	,
(	39192	)	,
(	39175	)	,
(	39158	)	,
(	39141	)	,
(	39124	)	,
(	39107	)	,
(	39090	)	,
(	39073	)	,
(	39056	)	,
(	39039	)	,
(	39022	)	,
(	39005	)	,
(	38988	)	,
(	38971	)	,
(	38954	)	,
(	38937	)	,
(	38920	)	,
(	38903	)	,
(	38886	)	,
(	38869	)	,
(	38852	)	,
(	38835	)	,
(	38818	)	,
(	38801	)	,
(	38784	)	,
(	38767	)	,
(	38750	)	,
(	38733	)	,
(	38716	)	,
(	38699	)	,
(	38682	)	,
(	38665	)	,
(	38648	)	,
(	38631	)	,
(	38614	)	,
(	38597	)	,
(	38580	)	,
(	38563	)	,
(	38546	)	,
(	38529	)	,
(	38512	)	,
(	38495	)	,
(	38478	)	,
(	38461	)	,
(	38444	)	,
(	38427	)	,
(	38410	)	,
(	38393	)	,
(	38376	)	,
(	38359	)	,
(	38342	)	,
(	38325	)	,
(	38308	)	,
(	38291	)	,
(	38274	)	,
(	38257	)	,
(	38240	)	,
(	38223	)	,
(	38206	)	,
(	38189	)	,
(	38172	)	,
(	38155	)	,
(	38138	)	,
(	38121	)	,
(	38104	)	,
(	38087	)	,
(	38070	)	,
(	38053	)	,
(	38036	)	,
(	38019	)	,
(	38002	)	,
(	37985	)	,
(	37968	)	,
(	37951	)	,
(	37934	)	,
(	37917	)	,
(	37900	)	,
(	37883	)	,
(	37866	)	,
(	37849	)	,
(	37832	)	,
(	37815	)	,
(	37798	)	,
(	37781	)	,
(	37764	)	,
(	37747	)	,
(	37730	)	,
(	37713	)	,
(	37696	)	,
(	37679	)	,
(	37662	)	,
(	37645	)	,
(	37628	)	,
(	37611	)	,
(	37594	)	,
(	37577	)	,
(	37560	)	,
(	37543	)	,
(	37526	)	,
(	37509	)	,
(	37492	)	,
(	37475	)	,
(	37458	)	,
(	37441	)	,
(	37424	)	,
(	37407	)	,
(	37390	)	,
(	37373	)	,
(	37356	)	,
(	37339	)	,
(	37322	)	,
(	37305	)	,
(	37288	)	,
(	37271	)	,
(	37254	)	,
(	37237	)	,
(	37220	)	,
(	37203	)	,
(	37186	)	,
(	37169	)	,
(	37152	)	,
(	37135	)	,
(	37118	)	,
(	37101	)	,
(	37084	)	,
(	37067	)	,
(	37050	)	,
(	37033	)	,
(	37016	)	,
(	36999	)	,
(	36982	)	,
(	36965	)	,
(	36948	)	,
(	36931	)	,
(	36914	)	,
(	36897	)	,
(	36880	)	,
(	36863	)	,
(	36846	)	,
(	36829	)	,
(	36812	)	,
(	36795	)	,
(	36778	)	,
(	36761	)	,
(	36744	)	,
(	36727	)	,
(	36710	)	,
(	36693	)	,
(	36676	)	,
(	36659	)	,
(	36642	)	,
(	36625	)	,
(	36608	)	,
(	36591	)	,
(	36574	)	,
(	36557	)	,
(	36540	)	,
(	36523	)	,
(	36506	)	,
(	36489	)	,
(	36472	)	,
(	36455	)	,
(	36438	)	,
(	36421	)	,
(	36404	)	,
(	36387	)	,
(	36370	)	,
(	36353	)	,
(	36336	)	,
(	36319	)	,
(	36302	)	,
(	36285	)	,
(	36268	)	,
(	36251	)	,
(	36234	)	,
(	36217	)	,
(	36200	)	,
(	36183	)	,
(	36166	)	,
(	36149	)	,
(	36132	)	,
(	36115	)	,
(	36098	)	,
(	36081	)	,
(	36064	)	,
(	36047	)	,
(	36030	)	,
(	36013	)	,
(	35996	)	,
(	35979	)	,
(	35962	)	,
(	35945	)	,
(	35928	)	,
(	35911	)	,
(	35894	)	,
(	35877	)	,
(	35860	)	,
(	35843	)	,
(	35826	)	,
(	35809	)	,
(	35792	)	,
(	35775	)	,
(	35758	)	,
(	35741	)	,
(	35724	)	,
(	35707	)	,
(	35690	)	,
(	35673	)	,
(	35656	)	,
(	35639	)	,
(	35622	)	,
(	35605	)	,
(	35588	)	,
(	35571	)	,
(	35554	)	,
(	35537	)	,
(	35520	)	,
(	35503	)	,
(	35486	)	,
(	35469	)	,
(	35452	)	,
(	35435	)	,
(	35418	)	,
(	35401	)	,
(	35384	)	,
(	35367	)	,
(	35350	)	,
(	35333	)	,
(	35316	)	,
(	35299	)	,
(	35282	)	,
(	35265	)	,
(	35248	)	,
(	35231	)	,
(	35214	)	,
(	35197	)	,
(	35180	)	,
(	35163	)	,
(	35146	)	,
(	35129	)	,
(	35112	)	,
(	35095	)	,
(	35078	)	,
(	35061	)	,
(	35044	)	,
(	35027	)	,
(	35010	)	,
(	34993	)	,
(	34976	)	,
(	34959	)	,
(	34942	)	,
(	34925	)	,
(	34908	)	,
(	34891	)	,
(	34874	)	,
(	34857	)	,
(	34840	)	,
(	34823	)	,
(	34806	)	,
(	34789	)	,
(	34772	)	,
(	34755	)	,
(	34738	)	,
(	34721	)	,
(	34704	)	,
(	34687	)	,
(	34670	)	,
(	34653	)	,
(	34636	)	,
(	34619	)	,
(	34602	)	,
(	34585	)	,
(	34568	)	,
(	34551	)	,
(	34534	)	,
(	34517	)	,
(	34500	)	,
(	34483	)	,
(	34466	)	,
(	34449	)	,
(	34432	)	,
(	34415	)	,
(	34398	)	,
(	34381	)	,
(	34364	)	,
(	34347	)	,
(	34330	)	,
(	34313	)	,
(	34296	)	,
(	34279	)	,
(	34262	)	,
(	34245	)	,
(	34228	)	,
(	34211	)	,
(	34194	)	,
(	34177	)	,
(	34160	)	,
(	34143	)	,
(	34126	)	,
(	34109	)	,
(	34092	)	,
(	34075	)	,
(	34058	)	,
(	34041	)	,
(	34024	)	,
(	34007	)	,
(	33990	)	,
(	33973	)	,
(	33956	)	,
(	33939	)	,
(	33922	)	,
(	33905	)	,
(	33888	)	,
(	33871	)	,
(	33854	)	,
(	33837	)	,
(	33820	)	,
(	33803	)	,
(	33786	)	,
(	33769	)	,
(	33752	)	,
(	33735	)	,
(	33718	)	,
(	33701	)	,
(	33684	)	,
(	33667	)	,
(	33650	)	,
(	33633	)	,
(	33616	)	,
(	33599	)	,
(	33582	)	,
(	33565	)	,
(	33548	)	,
(	33531	)	,
(	33514	)	,
(	33497	)	,
(	33480	)	,
(	33463	)	,
(	33446	)	,
(	33429	)	,
(	33412	)	,
(	33395	)	,
(	33378	)	,
(	33361	)	,
(	33344	)	,
(	33327	)	,
(	33310	)	,
(	33293	)	,
(	33276	)	,
(	33259	)	,
(	33242	)	,
(	33225	)	,
(	33208	)	,
(	33191	)	,
(	33174	)	,
(	33157	)	,
(	33140	)	,
(	33123	)	,
(	33106	)	,
(	33089	)	,
(	33072	)	,
(	33055	)	,
(	33038	)	,
(	33021	)	,
(	33004	)	,
(	32987	)	,
(	32970	)	,
(	32953	)	,
(	32936	)	,
(	32919	)	,
(	32902	)	,
(	32885	)	,
(	32868	)	,
(	32851	)	,
(	32834	)	,
(	32817	)	,
(	32800	)	,
(	32783	)	,
(	32766	)	,
(	32749	)	,
(	32732	)	,
(	32715	)	,
(	32698	)	,
(	32681	)	,
(	32664	)	,
(	32647	)	,
(	32630	)	,
(	32613	)	,
(	32596	)	,
(	32579	)	,
(	32562	)	,
(	32545	)	,
(	32528	)	,
(	32511	)	,
(	32494	)	,
(	32477	)	,
(	32460	)	,
(	32443	)	,
(	32426	)	,
(	32409	)	,
(	32392	)	,
(	32375	)	,
(	32358	)	,
(	32341	)	,
(	32324	)	,
(	32307	)	,
(	32290	)	,
(	32273	)	,
(	32256	)	,
(	32239	)	,
(	32222	)	,
(	32205	)	,
(	32188	)	,
(	32171	)	,
(	32154	)	,
(	32137	)	,
(	32120	)	,
(	32103	)	,
(	32086	)	,
(	32069	)	,
(	32052	)	,
(	32035	)	,
(	32018	)	,
(	32001	)	,
(	31984	)	,
(	31967	)	,
(	31950	)	,
(	31933	)	,
(	31916	)	,
(	31899	)	,
(	31882	)	,
(	31865	)	,
(	31848	)	,
(	31831	)	,
(	31814	)	,
(	31797	)	,
(	31780	)	,
(	31763	)	,
(	31746	)	,
(	31729	)	,
(	31712	)	,
(	31695	)	,
(	31678	)	,
(	31661	)	,
(	31644	)	,
(	31627	)	,
(	31610	)	,
(	31593	)	,
(	31576	)	,
(	31559	)	,
(	31542	)	,
(	31525	)	,
(	31508	)	,
(	31491	)	,
(	31474	)	,
(	31457	)	,
(	31440	)	,
(	31423	)	,
(	31406	)	,
(	31389	)	,
(	31372	)	,
(	31355	)	,
(	31338	)	,
(	31321	)	,
(	31304	)	,
(	31287	)	,
(	31270	)	,
(	31253	)	,
(	31236	)	,
(	31219	)	,
(	31202	)	,
(	31185	)	,
(	31168	)	,
(	31151	)	,
(	31134	)	,
(	31117	)	,
(	31100	)	,
(	31083	)	,
(	31066	)	,
(	31049	)	,
(	31032	)	,
(	31015	)	,
(	30998	)	,
(	30981	)	,
(	30964	)	,
(	30947	)	,
(	30930	)	,
(	30913	)	,
(	30896	)	,
(	30879	)	,
(	30862	)	,
(	30845	)	,
(	30828	)	,
(	30811	)	,
(	30794	)	,
(	30777	)	,
(	30760	)	,
(	30743	)	,
(	30726	)	,
(	30709	)	,
(	30692	)	,
(	30675	)	,
(	30658	)	,
(	30641	)	,
(	30624	)	,
(	30607	)	,
(	30590	)	,
(	30573	)	,
(	30556	)	,
(	30539	)	,
(	30522	)	,
(	30505	)	,
(	30488	)	,
(	30471	)	,
(	30454	)	,
(	30437	)	,
(	30420	)	,
(	30403	)	,
(	30386	)	,
(	30369	)	,
(	30352	)	,
(	30335	)	,
(	30318	)	,
(	30301	)	,
(	30284	)	,
(	30267	)	,
(	30250	)	,
(	30233	)	,
(	30216	)	,
(	30199	)	,
(	30182	)	,
(	30165	)	,
(	30148	)	,
(	30131	)	,
(	30114	)	,
(	30097	)	,
(	30080	)	,
(	30063	)	,
(	30046	)	,
(	30029	)	,
(	30012	)	,
(	29995	)	,
(	29978	)	,
(	29961	)	,
(	29944	)	,
(	29927	)	,
(	29910	)	,
(	29893	)	,
(	29876	)	,
(	29859	)	,
(	29842	)	,
(	29825	)	,
(	29808	)	,
(	29791	)	,
(	29774	)	,
(	29757	)	,
(	29740	)	,
(	29723	)	,
(	29706	)	,
(	29689	)	,
(	29672	)	,
(	29655	)	,
(	29638	)	,
(	29621	)	,
(	29604	)	,
(	29587	)	,
(	29570	)	,
(	29553	)	,
(	29536	)	,
(	29519	)	,
(	29502	)	,
(	29485	)	,
(	29468	)	,
(	29451	)	,
(	29434	)	,
(	29417	)	,
(	29400	)	,
(	29383	)	,
(	29366	)	,
(	29349	)	,
(	29332	)	,
(	29315	)	,
(	29298	)	,
(	29281	)	,
(	29264	)	,
(	29247	)	,
(	29230	)	,
(	29213	)	,
(	29196	)	,
(	29179	)	,
(	29162	)	,
(	29145	)	,
(	29128	)	,
(	29111	)	,
(	29094	)	,
(	29077	)	,
(	29060	)	,
(	29043	)	,
(	29026	)	,
(	29009	)	,
(	28992	)	,
(	28975	)	,
(	28958	)	,
(	28941	)	,
(	28924	)	,
(	28907	)	,
(	28890	)	,
(	28873	)	,
(	28856	)	,
(	28839	)	,
(	28822	)	,
(	28805	)	,
(	28788	)	,
(	28771	)	,
(	28754	)	,
(	28737	)	,
(	28720	)	,
(	28703	)	,
(	28686	)	,
(	28669	)	,
(	28652	)	,
(	28635	)	,
(	28618	)	,
(	28601	)	,
(	28584	)	,
(	28567	)	,
(	28550	)	,
(	28533	)	,
(	28516	)	,
(	28499	)	,
(	28482	)	,
(	28465	)	,
(	28448	)	,
(	28431	)	,
(	28414	)	,
(	28397	)	,
(	28380	)	,
(	28363	)	,
(	28346	)	,
(	28329	)	,
(	28312	)	,
(	28295	)	,
(	28278	)	,
(	28261	)	,
(	28244	)	,
(	28227	)	,
(	28210	)	,
(	28193	)	,
(	28176	)	,
(	28159	)	,
(	28142	)	,
(	28125	)	,
(	28108	)	,
(	28091	)	,
(	28074	)	,
(	28057	)	,
(	28040	)	,
(	28023	)	,
(	28006	)	,
(	27989	)	,
(	27972	)	,
(	27955	)	,
(	27938	)	,
(	27921	)	,
(	27904	)	,
(	27887	)	,
(	27870	)	,
(	27853	)	,
(	27836	)	,
(	27819	)	,
(	27802	)	,
(	27785	)	,
(	27768	)	,
(	27751	)	,
(	27734	)	,
(	27717	)	,
(	27700	)	,
(	27683	)	,
(	27666	)	,
(	27649	)	,
(	27632	)	,
(	27615	)	,
(	27598	)	,
(	27581	)	,
(	27564	)	,
(	27547	)	,
(	27530	)	,
(	27513	)	,
(	27496	)	,
(	27479	)	,
(	27462	)	,
(	27445	)	,
(	27428	)	,
(	27411	)	,
(	27394	)	,
(	27377	)	,
(	27360	)	,
(	27343	)	,
(	27326	)	,
(	27309	)	,
(	27292	)	,
(	27275	)	,
(	27258	)	,
(	27241	)	,
(	27224	)	,
(	27207	)	,
(	27190	)	,
(	27173	)	,
(	27156	)	,
(	27139	)	,
(	27122	)	,
(	27105	)	,
(	27088	)	,
(	27071	)	,
(	27054	)	,
(	27037	)	,
(	27020	)	,
(	27003	)	,
(	26986	)	,
(	26969	)	,
(	26952	)	,
(	26935	)	,
(	26918	)	,
(	26901	)	,
(	26884	)	,
(	26867	)	,
(	26850	)	,
(	26833	)	,
(	26816	)	,
(	26799	)	,
(	26782	)	,
(	26765	)	,
(	26748	)	,
(	26731	)	,
(	26714	)	,
(	26697	)	,
(	26680	)	,
(	26663	)	,
(	26646	)	,
(	26629	)	,
(	26612	)	,
(	26595	)	,
(	26578	)	,
(	26561	)	,
(	26544	)	,
(	26527	)	,
(	26510	)	,
(	26493	)	,
(	26476	)	,
(	26459	)	,
(	26442	)	,
(	26425	)	,
(	26408	)	,
(	26391	)	,
(	26374	)	,
(	26357	)	,
(	26340	)	,
(	26323	)	,
(	26306	)	,
(	26289	)	,
(	26272	)	,
(	26255	)	,
(	26238	)	,
(	26221	)	,
(	26204	)	,
(	26187	)	,
(	26170	)	,
(	26153	)	,
(	26136	)	,
(	26119	)	,
(	26102	)	,
(	26085	)	,
(	26068	)	,
(	26051	)	,
(	26034	)	,
(	26017	)	,
(	26000	)	

 );
 
 end package LED_Flash_LUT_pkg;