library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package buzzer_LUT_pkg is
 
 type my_array is array (4095 downto 0) of integer;
 constant DtoBP_LUT : my_array := ( -- can this be the same name as the one used for the display?
 
(	17500	)	,
(	17496	)	,
(	17492	)	,
(	17488	)	,
(	17484	)	,
(	17480	)	,
(	17476	)	,
(	17472	)	,
(	17468	)	,
(	17464	)	,
(	17460	)	,
(	17456	)	,
(	17452	)	,
(	17448	)	,
(	17444	)	,
(	17440	)	,
(	17436	)	,
(	17432	)	,
(	17428	)	,
(	17424	)	,
(	17420	)	,
(	17416	)	,
(	17412	)	,
(	17408	)	,
(	17404	)	,
(	17400	)	,
(	17396	)	,
(	17392	)	,
(	17388	)	,
(	17384	)	,
(	17380	)	,
(	17376	)	,
(	17372	)	,
(	17368	)	,
(	17364	)	,
(	17360	)	,
(	17356	)	,
(	17352	)	,
(	17348	)	,
(	17344	)	,
(	17340	)	,
(	17336	)	,
(	17332	)	,
(	17328	)	,
(	17324	)	,
(	17320	)	,
(	17316	)	,
(	17312	)	,
(	17308	)	,
(	17304	)	,
(	17300	)	,
(	17296	)	,
(	17292	)	,
(	17288	)	,
(	17284	)	,
(	17280	)	,
(	17276	)	,
(	17272	)	,
(	17268	)	,
(	17264	)	,
(	17260	)	,
(	17256	)	,
(	17252	)	,
(	17248	)	,
(	17244	)	,
(	17240	)	,
(	17236	)	,
(	17232	)	,
(	17228	)	,
(	17224	)	,
(	17220	)	,
(	17216	)	,
(	17212	)	,
(	17208	)	,
(	17204	)	,
(	17200	)	,
(	17196	)	,
(	17192	)	,
(	17188	)	,
(	17184	)	,
(	17180	)	,
(	17176	)	,
(	17172	)	,
(	17168	)	,
(	17164	)	,
(	17160	)	,
(	17156	)	,
(	17152	)	,
(	17148	)	,
(	17144	)	,
(	17140	)	,
(	17136	)	,
(	17132	)	,
(	17128	)	,
(	17124	)	,
(	17120	)	,
(	17116	)	,
(	17112	)	,
(	17108	)	,
(	17104	)	,
(	17100	)	,
(	17096	)	,
(	17092	)	,
(	17088	)	,
(	17084	)	,
(	17080	)	,
(	17076	)	,
(	17072	)	,
(	17068	)	,
(	17064	)	,
(	17060	)	,
(	17056	)	,
(	17052	)	,
(	17048	)	,
(	17044	)	,
(	17040	)	,
(	17036	)	,
(	17032	)	,
(	17028	)	,
(	17024	)	,
(	17020	)	,
(	17016	)	,
(	17012	)	,
(	17008	)	,
(	17004	)	,
(	17000	)	,
(	16996	)	,
(	16992	)	,
(	16988	)	,
(	16984	)	,
(	16980	)	,
(	16976	)	,
(	16972	)	,
(	16968	)	,
(	16964	)	,
(	16960	)	,
(	16956	)	,
(	16952	)	,
(	16948	)	,
(	16944	)	,
(	16940	)	,
(	16936	)	,
(	16932	)	,
(	16928	)	,
(	16924	)	,
(	16920	)	,
(	16916	)	,
(	16912	)	,
(	16908	)	,
(	16904	)	,
(	16900	)	,
(	16896	)	,
(	16892	)	,
(	16888	)	,
(	16884	)	,
(	16880	)	,
(	16876	)	,
(	16872	)	,
(	16868	)	,
(	16864	)	,
(	16860	)	,
(	16856	)	,
(	16852	)	,
(	16848	)	,
(	16844	)	,
(	16840	)	,
(	16836	)	,
(	16832	)	,
(	16828	)	,
(	16824	)	,
(	16820	)	,
(	16816	)	,
(	16812	)	,
(	16808	)	,
(	16804	)	,
(	16800	)	,
(	16796	)	,
(	16792	)	,
(	16788	)	,
(	16784	)	,
(	16780	)	,
(	16776	)	,
(	16772	)	,
(	16768	)	,
(	16764	)	,
(	16760	)	,
(	16756	)	,
(	16752	)	,
(	16748	)	,
(	16744	)	,
(	16740	)	,
(	16736	)	,
(	16732	)	,
(	16728	)	,
(	16724	)	,
(	16720	)	,
(	16716	)	,
(	16712	)	,
(	16708	)	,
(	16704	)	,
(	16700	)	,
(	16696	)	,
(	16692	)	,
(	16688	)	,
(	16684	)	,
(	16680	)	,
(	16676	)	,
(	16672	)	,
(	16668	)	,
(	16664	)	,
(	16660	)	,
(	16656	)	,
(	16652	)	,
(	16648	)	,
(	16644	)	,
(	16640	)	,
(	16636	)	,
(	16632	)	,
(	16628	)	,
(	16624	)	,
(	16620	)	,
(	16616	)	,
(	16612	)	,
(	16608	)	,
(	16604	)	,
(	16600	)	,
(	16596	)	,
(	16592	)	,
(	16588	)	,
(	16584	)	,
(	16580	)	,
(	16576	)	,
(	16572	)	,
(	16568	)	,
(	16564	)	,
(	16560	)	,
(	16556	)	,
(	16552	)	,
(	16548	)	,
(	16544	)	,
(	16540	)	,
(	16536	)	,
(	16532	)	,
(	16528	)	,
(	16524	)	,
(	16520	)	,
(	16516	)	,
(	16512	)	,
(	16508	)	,
(	16504	)	,
(	16500	)	,
(	16496	)	,
(	16492	)	,
(	16488	)	,
(	16484	)	,
(	16480	)	,
(	16476	)	,
(	16472	)	,
(	16468	)	,
(	16464	)	,
(	16460	)	,
(	16456	)	,
(	16452	)	,
(	16448	)	,
(	16444	)	,
(	16440	)	,
(	16436	)	,
(	16432	)	,
(	16428	)	,
(	16424	)	,
(	16420	)	,
(	16416	)	,
(	16412	)	,
(	16408	)	,
(	16404	)	,
(	16400	)	,
(	16396	)	,
(	16392	)	,
(	16388	)	,
(	16384	)	,
(	16380	)	,
(	16376	)	,
(	16372	)	,
(	16368	)	,
(	16364	)	,
(	16360	)	,
(	16356	)	,
(	16352	)	,
(	16348	)	,
(	16344	)	,
(	16340	)	,
(	16336	)	,
(	16332	)	,
(	16328	)	,
(	16324	)	,
(	16320	)	,
(	16316	)	,
(	16312	)	,
(	16308	)	,
(	16304	)	,
(	16300	)	,
(	16296	)	,
(	16292	)	,
(	16288	)	,
(	16284	)	,
(	16280	)	,
(	16276	)	,
(	16272	)	,
(	16268	)	,
(	16264	)	,
(	16260	)	,
(	16256	)	,
(	16252	)	,
(	16248	)	,
(	16244	)	,
(	16240	)	,
(	16236	)	,
(	16232	)	,
(	16228	)	,
(	16224	)	,
(	16220	)	,
(	16216	)	,
(	16212	)	,
(	16208	)	,
(	16204	)	,
(	16200	)	,
(	16196	)	,
(	16192	)	,
(	16188	)	,
(	16184	)	,
(	16180	)	,
(	16176	)	,
(	16172	)	,
(	16168	)	,
(	16164	)	,
(	16160	)	,
(	16156	)	,
(	16152	)	,
(	16148	)	,
(	16144	)	,
(	16140	)	,
(	16136	)	,
(	16132	)	,
(	16128	)	,
(	16124	)	,
(	16120	)	,
(	16116	)	,
(	16112	)	,
(	16108	)	,
(	16104	)	,
(	16100	)	,
(	16096	)	,
(	16092	)	,
(	16088	)	,
(	16084	)	,
(	16080	)	,
(	16076	)	,
(	16072	)	,
(	16068	)	,
(	16064	)	,
(	16060	)	,
(	16056	)	,
(	16052	)	,
(	16048	)	,
(	16044	)	,
(	16040	)	,
(	16036	)	,
(	16032	)	,
(	16028	)	,
(	16024	)	,
(	16020	)	,
(	16016	)	,
(	16012	)	,
(	16008	)	,
(	16004	)	,
(	16000	)	,
(	15996	)	,
(	15992	)	,
(	15988	)	,
(	15984	)	,
(	15980	)	,
(	15976	)	,
(	15972	)	,
(	15968	)	,
(	15964	)	,
(	15960	)	,
(	15956	)	,
(	15952	)	,
(	15948	)	,
(	15944	)	,
(	15940	)	,
(	15936	)	,
(	15932	)	,
(	15928	)	,
(	15924	)	,
(	15920	)	,
(	15916	)	,
(	15912	)	,
(	15908	)	,
(	15904	)	,
(	15900	)	,
(	15896	)	,
(	15892	)	,
(	15888	)	,
(	15884	)	,
(	15880	)	,
(	15876	)	,
(	15872	)	,
(	15868	)	,
(	15864	)	,
(	15860	)	,
(	15856	)	,
(	15852	)	,
(	15848	)	,
(	15844	)	,
(	15840	)	,
(	15836	)	,
(	15832	)	,
(	15828	)	,
(	15824	)	,
(	15820	)	,
(	15816	)	,
(	15812	)	,
(	15808	)	,
(	15804	)	,
(	15800	)	,
(	15796	)	,
(	15792	)	,
(	15788	)	,
(	15784	)	,
(	15780	)	,
(	15776	)	,
(	15772	)	,
(	15768	)	,
(	15764	)	,
(	15760	)	,
(	15756	)	,
(	15752	)	,
(	15748	)	,
(	15744	)	,
(	15740	)	,
(	15736	)	,
(	15732	)	,
(	15728	)	,
(	15724	)	,
(	15720	)	,
(	15716	)	,
(	15712	)	,
(	15708	)	,
(	15704	)	,
(	15700	)	,
(	15696	)	,
(	15692	)	,
(	15688	)	,
(	15684	)	,
(	15680	)	,
(	15676	)	,
(	15672	)	,
(	15668	)	,
(	15664	)	,
(	15660	)	,
(	15656	)	,
(	15652	)	,
(	15648	)	,
(	15644	)	,
(	15640	)	,
(	15636	)	,
(	15632	)	,
(	15628	)	,
(	15624	)	,
(	15620	)	,
(	15616	)	,
(	15612	)	,
(	15608	)	,
(	15604	)	,
(	15600	)	,
(	15596	)	,
(	15592	)	,
(	15588	)	,
(	15584	)	,
(	15580	)	,
(	15576	)	,
(	15572	)	,
(	15568	)	,
(	15564	)	,
(	15560	)	,
(	15556	)	,
(	15552	)	,
(	15548	)	,
(	15544	)	,
(	15540	)	,
(	15536	)	,
(	15532	)	,
(	15528	)	,
(	15524	)	,
(	15520	)	,
(	15516	)	,
(	15512	)	,
(	15508	)	,
(	15504	)	,
(	15500	)	,
(	15496	)	,
(	15492	)	,
(	15488	)	,
(	15484	)	,
(	15480	)	,
(	15476	)	,
(	15472	)	,
(	15468	)	,
(	15464	)	,
(	15460	)	,
(	15456	)	,
(	15452	)	,
(	15448	)	,
(	15444	)	,
(	15440	)	,
(	15436	)	,
(	15432	)	,
(	15428	)	,
(	15424	)	,
(	15420	)	,
(	15416	)	,
(	15412	)	,
(	15408	)	,
(	15404	)	,
(	15400	)	,
(	15396	)	,
(	15392	)	,
(	15388	)	,
(	15384	)	,
(	15380	)	,
(	15376	)	,
(	15372	)	,
(	15368	)	,
(	15364	)	,
(	15360	)	,
(	15356	)	,
(	15352	)	,
(	15348	)	,
(	15344	)	,
(	15340	)	,
(	15336	)	,
(	15332	)	,
(	15328	)	,
(	15324	)	,
(	15320	)	,
(	15316	)	,
(	15312	)	,
(	15308	)	,
(	15304	)	,
(	15300	)	,
(	15296	)	,
(	15292	)	,
(	15288	)	,
(	15284	)	,
(	15280	)	,
(	15276	)	,
(	15272	)	,
(	15268	)	,
(	15264	)	,
(	15260	)	,
(	15256	)	,
(	15252	)	,
(	15248	)	,
(	15244	)	,
(	15240	)	,
(	15236	)	,
(	15232	)	,
(	15228	)	,
(	15224	)	,
(	15220	)	,
(	15216	)	,
(	15212	)	,
(	15208	)	,
(	15204	)	,
(	15200	)	,
(	15196	)	,
(	15192	)	,
(	15188	)	,
(	15184	)	,
(	15180	)	,
(	15176	)	,
(	15172	)	,
(	15168	)	,
(	15164	)	,
(	15160	)	,
(	15156	)	,
(	15152	)	,
(	15148	)	,
(	15144	)	,
(	15140	)	,
(	15136	)	,
(	15132	)	,
(	15128	)	,
(	15124	)	,
(	15120	)	,
(	15116	)	,
(	15112	)	,
(	15108	)	,
(	15104	)	,
(	15100	)	,
(	15096	)	,
(	15092	)	,
(	15088	)	,
(	15084	)	,
(	15080	)	,
(	15076	)	,
(	15072	)	,
(	15068	)	,
(	15064	)	,
(	15060	)	,
(	15056	)	,
(	15052	)	,
(	15048	)	,
(	15044	)	,
(	15040	)	,
(	15036	)	,
(	15032	)	,
(	15028	)	,
(	15024	)	,
(	15020	)	,
(	15016	)	,
(	15012	)	,
(	15008	)	,
(	15004	)	,
(	15000	)	,
(	14996	)	,
(	14992	)	,
(	14988	)	,
(	14984	)	,
(	14980	)	,
(	14976	)	,
(	14972	)	,
(	14968	)	,
(	14964	)	,
(	14960	)	,
(	14956	)	,
(	14952	)	,
(	14948	)	,
(	14944	)	,
(	14940	)	,
(	14936	)	,
(	14932	)	,
(	14928	)	,
(	14924	)	,
(	14920	)	,
(	14916	)	,
(	14912	)	,
(	14908	)	,
(	14904	)	,
(	14900	)	,
(	14896	)	,
(	14892	)	,
(	14888	)	,
(	14884	)	,
(	14880	)	,
(	14876	)	,
(	14872	)	,
(	14868	)	,
(	14864	)	,
(	14860	)	,
(	14856	)	,
(	14852	)	,
(	14848	)	,
(	14844	)	,
(	14840	)	,
(	14836	)	,
(	14832	)	,
(	14828	)	,
(	14824	)	,
(	14820	)	,
(	14816	)	,
(	14812	)	,
(	14808	)	,
(	14804	)	,
(	14800	)	,
(	14796	)	,
(	14792	)	,
(	14788	)	,
(	14784	)	,
(	14780	)	,
(	14776	)	,
(	14772	)	,
(	14768	)	,
(	14764	)	,
(	14760	)	,
(	14756	)	,
(	14752	)	,
(	14748	)	,
(	14744	)	,
(	14740	)	,
(	14736	)	,
(	14732	)	,
(	14728	)	,
(	14724	)	,
(	14720	)	,
(	14716	)	,
(	14712	)	,
(	14708	)	,
(	14704	)	,
(	14700	)	,
(	14696	)	,
(	14692	)	,
(	14688	)	,
(	14684	)	,
(	14680	)	,
(	14676	)	,
(	14672	)	,
(	14668	)	,
(	14664	)	,
(	14660	)	,
(	14656	)	,
(	14652	)	,
(	14648	)	,
(	14644	)	,
(	14640	)	,
(	14636	)	,
(	14632	)	,
(	14628	)	,
(	14624	)	,
(	14620	)	,
(	14616	)	,
(	14612	)	,
(	14608	)	,
(	14604	)	,
(	14600	)	,
(	14596	)	,
(	14592	)	,
(	14588	)	,
(	14584	)	,
(	14580	)	,
(	14576	)	,
(	14572	)	,
(	14568	)	,
(	14564	)	,
(	14560	)	,
(	14556	)	,
(	14552	)	,
(	14548	)	,
(	14544	)	,
(	14540	)	,
(	14536	)	,
(	14532	)	,
(	14528	)	,
(	14524	)	,
(	14520	)	,
(	14516	)	,
(	14512	)	,
(	14508	)	,
(	14504	)	,
(	14500	)	,
(	14496	)	,
(	14492	)	,
(	14488	)	,
(	14484	)	,
(	14480	)	,
(	14476	)	,
(	14472	)	,
(	14468	)	,
(	14464	)	,
(	14460	)	,
(	14456	)	,
(	14452	)	,
(	14448	)	,
(	14444	)	,
(	14440	)	,
(	14436	)	,
(	14432	)	,
(	14428	)	,
(	14424	)	,
(	14420	)	,
(	14416	)	,
(	14412	)	,
(	14408	)	,
(	14404	)	,
(	14400	)	,
(	14396	)	,
(	14392	)	,
(	14388	)	,
(	14384	)	,
(	14380	)	,
(	14376	)	,
(	14372	)	,
(	14368	)	,
(	14364	)	,
(	14360	)	,
(	14356	)	,
(	14352	)	,
(	14348	)	,
(	14344	)	,
(	14340	)	,
(	14336	)	,
(	14332	)	,
(	14328	)	,
(	14324	)	,
(	14320	)	,
(	14316	)	,
(	14312	)	,
(	14308	)	,
(	14304	)	,
(	14300	)	,
(	14296	)	,
(	14292	)	,
(	14288	)	,
(	14284	)	,
(	14280	)	,
(	14276	)	,
(	14272	)	,
(	14268	)	,
(	14264	)	,
(	14260	)	,
(	14256	)	,
(	14252	)	,
(	14248	)	,
(	14244	)	,
(	14240	)	,
(	14236	)	,
(	14232	)	,
(	14228	)	,
(	14224	)	,
(	14220	)	,
(	14216	)	,
(	14212	)	,
(	14208	)	,
(	14204	)	,
(	14200	)	,
(	14196	)	,
(	14192	)	,
(	14188	)	,
(	14184	)	,
(	14180	)	,
(	14176	)	,
(	14172	)	,
(	14168	)	,
(	14164	)	,
(	14160	)	,
(	14156	)	,
(	14152	)	,
(	14148	)	,
(	14144	)	,
(	14140	)	,
(	14136	)	,
(	14132	)	,
(	14128	)	,
(	14124	)	,
(	14120	)	,
(	14116	)	,
(	14112	)	,
(	14108	)	,
(	14104	)	,
(	14100	)	,
(	14096	)	,
(	14092	)	,
(	14088	)	,
(	14084	)	,
(	14080	)	,
(	14076	)	,
(	14072	)	,
(	14068	)	,
(	14064	)	,
(	14060	)	,
(	14056	)	,
(	14052	)	,
(	14048	)	,
(	14044	)	,
(	14040	)	,
(	14036	)	,
(	14032	)	,
(	14028	)	,
(	14024	)	,
(	14020	)	,
(	14016	)	,
(	14012	)	,
(	14008	)	,
(	14004	)	,
(	14000	)	,
(	13996	)	,
(	13992	)	,
(	13988	)	,
(	13984	)	,
(	13980	)	,
(	13976	)	,
(	13972	)	,
(	13968	)	,
(	13964	)	,
(	13960	)	,
(	13956	)	,
(	13952	)	,
(	13948	)	,
(	13944	)	,
(	13940	)	,
(	13936	)	,
(	13932	)	,
(	13928	)	,
(	13924	)	,
(	13920	)	,
(	13916	)	,
(	13912	)	,
(	13908	)	,
(	13904	)	,
(	13900	)	,
(	13896	)	,
(	13892	)	,
(	13888	)	,
(	13884	)	,
(	13880	)	,
(	13876	)	,
(	13872	)	,
(	13868	)	,
(	13864	)	,
(	13860	)	,
(	13856	)	,
(	13852	)	,
(	13848	)	,
(	13844	)	,
(	13840	)	,
(	13836	)	,
(	13832	)	,
(	13828	)	,
(	13824	)	,
(	13820	)	,
(	13816	)	,
(	13812	)	,
(	13808	)	,
(	13804	)	,
(	13800	)	,
(	13796	)	,
(	13792	)	,
(	13788	)	,
(	13784	)	,
(	13780	)	,
(	13776	)	,
(	13772	)	,
(	13768	)	,
(	13764	)	,
(	13760	)	,
(	13756	)	,
(	13752	)	,
(	13748	)	,
(	13744	)	,
(	13740	)	,
(	13736	)	,
(	13732	)	,
(	13728	)	,
(	13724	)	,
(	13720	)	,
(	13716	)	,
(	13712	)	,
(	13708	)	,
(	13704	)	,
(	13700	)	,
(	13696	)	,
(	13692	)	,
(	13688	)	,
(	13684	)	,
(	13680	)	,
(	13676	)	,
(	13672	)	,
(	13668	)	,
(	13664	)	,
(	13660	)	,
(	13656	)	,
(	13652	)	,
(	13648	)	,
(	13644	)	,
(	13640	)	,
(	13636	)	,
(	13632	)	,
(	13628	)	,
(	13624	)	,
(	13620	)	,
(	13616	)	,
(	13612	)	,
(	13608	)	,
(	13604	)	,
(	13600	)	,
(	13596	)	,
(	13592	)	,
(	13588	)	,
(	13584	)	,
(	13580	)	,
(	13576	)	,
(	13572	)	,
(	13568	)	,
(	13564	)	,
(	13560	)	,
(	13556	)	,
(	13552	)	,
(	13548	)	,
(	13544	)	,
(	13540	)	,
(	13536	)	,
(	13532	)	,
(	13528	)	,
(	13524	)	,
(	13520	)	,
(	13516	)	,
(	13512	)	,
(	13508	)	,
(	13504	)	,
(	13500	)	,
(	13496	)	,
(	13492	)	,
(	13488	)	,
(	13484	)	,
(	13480	)	,
(	13476	)	,
(	13472	)	,
(	13468	)	,
(	13464	)	,
(	13460	)	,
(	13456	)	,
(	13452	)	,
(	13448	)	,
(	13444	)	,
(	13440	)	,
(	13436	)	,
(	13432	)	,
(	13428	)	,
(	13424	)	,
(	13420	)	,
(	13416	)	,
(	13412	)	,
(	13408	)	,
(	13404	)	,
(	13400	)	,
(	13396	)	,
(	13392	)	,
(	13388	)	,
(	13384	)	,
(	13380	)	,
(	13376	)	,
(	13372	)	,
(	13368	)	,
(	13364	)	,
(	13360	)	,
(	13356	)	,
(	13352	)	,
(	13348	)	,
(	13344	)	,
(	13340	)	,
(	13336	)	,
(	13332	)	,
(	13328	)	,
(	13324	)	,
(	13320	)	,
(	13316	)	,
(	13312	)	,
(	13308	)	,
(	13304	)	,
(	13300	)	,
(	13296	)	,
(	13292	)	,
(	13288	)	,
(	13284	)	,
(	13280	)	,
(	13276	)	,
(	13272	)	,
(	13268	)	,
(	13264	)	,
(	13260	)	,
(	13256	)	,
(	13252	)	,
(	13248	)	,
(	13244	)	,
(	13240	)	,
(	13236	)	,
(	13232	)	,
(	13228	)	,
(	13224	)	,
(	13220	)	,
(	13216	)	,
(	13212	)	,
(	13208	)	,
(	13204	)	,
(	13200	)	,
(	13196	)	,
(	13192	)	,
(	13188	)	,
(	13184	)	,
(	13180	)	,
(	13176	)	,
(	13172	)	,
(	13168	)	,
(	13164	)	,
(	13160	)	,
(	13156	)	,
(	13152	)	,
(	13148	)	,
(	13144	)	,
(	13140	)	,
(	13136	)	,
(	13132	)	,
(	13128	)	,
(	13124	)	,
(	13120	)	,
(	13116	)	,
(	13112	)	,
(	13108	)	,
(	13104	)	,
(	13100	)	,
(	13096	)	,
(	13092	)	,
(	13088	)	,
(	13084	)	,
(	13080	)	,
(	13076	)	,
(	13072	)	,
(	13068	)	,
(	13064	)	,
(	13060	)	,
(	13056	)	,
(	13052	)	,
(	13048	)	,
(	13044	)	,
(	13040	)	,
(	13036	)	,
(	13032	)	,
(	13028	)	,
(	13024	)	,
(	13020	)	,
(	13016	)	,
(	13012	)	,
(	13008	)	,
(	13004	)	,
(	13000	)	,
(	12996	)	,
(	12992	)	,
(	12988	)	,
(	12984	)	,
(	12980	)	,
(	12976	)	,
(	12972	)	,
(	12968	)	,
(	12964	)	,
(	12960	)	,
(	12956	)	,
(	12952	)	,
(	12948	)	,
(	12944	)	,
(	12940	)	,
(	12936	)	,
(	12932	)	,
(	12928	)	,
(	12924	)	,
(	12920	)	,
(	12916	)	,
(	12912	)	,
(	12908	)	,
(	12904	)	,
(	12900	)	,
(	12896	)	,
(	12892	)	,
(	12888	)	,
(	12884	)	,
(	12880	)	,
(	12876	)	,
(	12872	)	,
(	12868	)	,
(	12864	)	,
(	12860	)	,
(	12856	)	,
(	12852	)	,
(	12848	)	,
(	12844	)	,
(	12840	)	,
(	12836	)	,
(	12832	)	,
(	12828	)	,
(	12824	)	,
(	12820	)	,
(	12816	)	,
(	12812	)	,
(	12808	)	,
(	12804	)	,
(	12800	)	,
(	12796	)	,
(	12792	)	,
(	12788	)	,
(	12784	)	,
(	12780	)	,
(	12776	)	,
(	12772	)	,
(	12768	)	,
(	12764	)	,
(	12760	)	,
(	12756	)	,
(	12752	)	,
(	12748	)	,
(	12744	)	,
(	12740	)	,
(	12736	)	,
(	12732	)	,
(	12728	)	,
(	12724	)	,
(	12720	)	,
(	12716	)	,
(	12712	)	,
(	12708	)	,
(	12704	)	,
(	12700	)	,
(	12696	)	,
(	12692	)	,
(	12688	)	,
(	12684	)	,
(	12680	)	,
(	12676	)	,
(	12672	)	,
(	12668	)	,
(	12664	)	,
(	12660	)	,
(	12656	)	,
(	12652	)	,
(	12648	)	,
(	12644	)	,
(	12640	)	,
(	12636	)	,
(	12632	)	,
(	12628	)	,
(	12624	)	,
(	12620	)	,
(	12616	)	,
(	12612	)	,
(	12608	)	,
(	12604	)	,
(	12600	)	,
(	12596	)	,
(	12592	)	,
(	12588	)	,
(	12584	)	,
(	12580	)	,
(	12576	)	,
(	12572	)	,
(	12568	)	,
(	12564	)	,
(	12560	)	,
(	12556	)	,
(	12552	)	,
(	12548	)	,
(	12544	)	,
(	12540	)	,
(	12536	)	,
(	12532	)	,
(	12528	)	,
(	12524	)	,
(	12520	)	,
(	12516	)	,
(	12512	)	,
(	12508	)	,
(	12504	)	,
(	12500	)	,
(	12496	)	,
(	12492	)	,
(	12488	)	,
(	12484	)	,
(	12480	)	,
(	12476	)	,
(	12472	)	,
(	12468	)	,
(	12464	)	,
(	12460	)	,
(	12456	)	,
(	12452	)	,
(	12448	)	,
(	12444	)	,
(	12440	)	,
(	12436	)	,
(	12432	)	,
(	12428	)	,
(	12424	)	,
(	12420	)	,
(	12416	)	,
(	12412	)	,
(	12408	)	,
(	12404	)	,
(	12400	)	,
(	12396	)	,
(	12392	)	,
(	12388	)	,
(	12384	)	,
(	12380	)	,
(	12376	)	,
(	12372	)	,
(	12368	)	,
(	12364	)	,
(	12360	)	,
(	12356	)	,
(	12352	)	,
(	12348	)	,
(	12344	)	,
(	12340	)	,
(	12336	)	,
(	12332	)	,
(	12328	)	,
(	12324	)	,
(	12320	)	,
(	12316	)	,
(	12312	)	,
(	12308	)	,
(	12304	)	,
(	12300	)	,
(	12296	)	,
(	12292	)	,
(	12288	)	,
(	12284	)	,
(	12280	)	,
(	12276	)	,
(	12272	)	,
(	12268	)	,
(	12264	)	,
(	12260	)	,
(	12256	)	,
(	12252	)	,
(	12248	)	,
(	12244	)	,
(	12240	)	,
(	12236	)	,
(	12232	)	,
(	12228	)	,
(	12224	)	,
(	12220	)	,
(	12216	)	,
(	12212	)	,
(	12208	)	,
(	12204	)	,
(	12200	)	,
(	12196	)	,
(	12192	)	,
(	12188	)	,
(	12184	)	,
(	12180	)	,
(	12176	)	,
(	12172	)	,
(	12168	)	,
(	12164	)	,
(	12160	)	,
(	12156	)	,
(	12152	)	,
(	12148	)	,
(	12144	)	,
(	12140	)	,
(	12136	)	,
(	12132	)	,
(	12128	)	,
(	12124	)	,
(	12120	)	,
(	12116	)	,
(	12112	)	,
(	12108	)	,
(	12104	)	,
(	12100	)	,
(	12096	)	,
(	12092	)	,
(	12088	)	,
(	12084	)	,
(	12080	)	,
(	12076	)	,
(	12072	)	,
(	12068	)	,
(	12064	)	,
(	12060	)	,
(	12056	)	,
(	12052	)	,
(	12048	)	,
(	12044	)	,
(	12040	)	,
(	12036	)	,
(	12032	)	,
(	12028	)	,
(	12024	)	,
(	12020	)	,
(	12016	)	,
(	12012	)	,
(	12008	)	,
(	12004	)	,
(	12000	)	,
(	11996	)	,
(	11992	)	,
(	11988	)	,
(	11984	)	,
(	11980	)	,
(	11976	)	,
(	11972	)	,
(	11968	)	,
(	11964	)	,
(	11960	)	,
(	11956	)	,
(	11952	)	,
(	11948	)	,
(	11944	)	,
(	11940	)	,
(	11936	)	,
(	11932	)	,
(	11928	)	,
(	11924	)	,
(	11920	)	,
(	11916	)	,
(	11912	)	,
(	11908	)	,
(	11904	)	,
(	11900	)	,
(	11896	)	,
(	11892	)	,
(	11888	)	,
(	11884	)	,
(	11880	)	,
(	11876	)	,
(	11872	)	,
(	11868	)	,
(	11864	)	,
(	11860	)	,
(	11856	)	,
(	11852	)	,
(	11848	)	,
(	11844	)	,
(	11840	)	,
(	11836	)	,
(	11832	)	,
(	11828	)	,
(	11824	)	,
(	11820	)	,
(	11816	)	,
(	11812	)	,
(	11808	)	,
(	11804	)	,
(	11800	)	,
(	11796	)	,
(	11792	)	,
(	11788	)	,
(	11784	)	,
(	11780	)	,
(	11776	)	,
(	11772	)	,
(	11768	)	,
(	11764	)	,
(	11760	)	,
(	11756	)	,
(	11752	)	,
(	11748	)	,
(	11744	)	,
(	11740	)	,
(	11736	)	,
(	11732	)	,
(	11728	)	,
(	11724	)	,
(	11720	)	,
(	11716	)	,
(	11712	)	,
(	11708	)	,
(	11704	)	,
(	11700	)	,
(	11696	)	,
(	11692	)	,
(	11688	)	,
(	11684	)	,
(	11680	)	,
(	11676	)	,
(	11672	)	,
(	11668	)	,
(	11664	)	,
(	11660	)	,
(	11656	)	,
(	11652	)	,
(	11648	)	,
(	11644	)	,
(	11640	)	,
(	11636	)	,
(	11632	)	,
(	11628	)	,
(	11624	)	,
(	11620	)	,
(	11616	)	,
(	11612	)	,
(	11608	)	,
(	11604	)	,
(	11600	)	,
(	11596	)	,
(	11592	)	,
(	11588	)	,
(	11584	)	,
(	11580	)	,
(	11576	)	,
(	11572	)	,
(	11568	)	,
(	11564	)	,
(	11560	)	,
(	11556	)	,
(	11552	)	,
(	11548	)	,
(	11544	)	,
(	11540	)	,
(	11536	)	,
(	11532	)	,
(	11528	)	,
(	11524	)	,
(	11520	)	,
(	11516	)	,
(	11512	)	,
(	11508	)	,
(	11504	)	,
(	11500	)	,
(	11496	)	,
(	11492	)	,
(	11488	)	,
(	11484	)	,
(	11480	)	,
(	11476	)	,
(	11472	)	,
(	11468	)	,
(	11464	)	,
(	11460	)	,
(	11456	)	,
(	11452	)	,
(	11448	)	,
(	11444	)	,
(	11440	)	,
(	11436	)	,
(	11432	)	,
(	11428	)	,
(	11424	)	,
(	11420	)	,
(	11416	)	,
(	11412	)	,
(	11408	)	,
(	11404	)	,
(	11400	)	,
(	11396	)	,
(	11392	)	,
(	11388	)	,
(	11384	)	,
(	11380	)	,
(	11376	)	,
(	11372	)	,
(	11368	)	,
(	11364	)	,
(	11360	)	,
(	11356	)	,
(	11352	)	,
(	11348	)	,
(	11344	)	,
(	11340	)	,
(	11336	)	,
(	11332	)	,
(	11328	)	,
(	11324	)	,
(	11320	)	,
(	11316	)	,
(	11312	)	,
(	11308	)	,
(	11304	)	,
(	11300	)	,
(	11296	)	,
(	11292	)	,
(	11288	)	,
(	11284	)	,
(	11280	)	,
(	11276	)	,
(	11272	)	,
(	11268	)	,
(	11264	)	,
(	11260	)	,
(	11256	)	,
(	11252	)	,
(	11248	)	,
(	11244	)	,
(	11240	)	,
(	11236	)	,
(	11232	)	,
(	11228	)	,
(	11224	)	,
(	11220	)	,
(	11216	)	,
(	11212	)	,
(	11208	)	,
(	11204	)	,
(	11200	)	,
(	11196	)	,
(	11192	)	,
(	11188	)	,
(	11184	)	,
(	11180	)	,
(	11176	)	,
(	11172	)	,
(	11168	)	,
(	11164	)	,
(	11160	)	,
(	11156	)	,
(	11152	)	,
(	11148	)	,
(	11144	)	,
(	11140	)	,
(	11136	)	,
(	11132	)	,
(	11128	)	,
(	11124	)	,
(	11120	)	,
(	11116	)	,
(	11112	)	,
(	11108	)	,
(	11104	)	,
(	11100	)	,
(	11096	)	,
(	11092	)	,
(	11088	)	,
(	11084	)	,
(	11080	)	,
(	11076	)	,
(	11072	)	,
(	11068	)	,
(	11064	)	,
(	11060	)	,
(	11056	)	,
(	11052	)	,
(	11048	)	,
(	11044	)	,
(	11040	)	,
(	11036	)	,
(	11032	)	,
(	11028	)	,
(	11024	)	,
(	11020	)	,
(	11016	)	,
(	11012	)	,
(	11008	)	,
(	11004	)	,
(	11000	)	,
(	10996	)	,
(	10992	)	,
(	10988	)	,
(	10984	)	,
(	10980	)	,
(	10976	)	,
(	10972	)	,
(	10968	)	,
(	10964	)	,
(	10960	)	,
(	10956	)	,
(	10952	)	,
(	10948	)	,
(	10944	)	,
(	10940	)	,
(	10936	)	,
(	10932	)	,
(	10928	)	,
(	10924	)	,
(	10920	)	,
(	10916	)	,
(	10912	)	,
(	10908	)	,
(	10904	)	,
(	10900	)	,
(	10896	)	,
(	10892	)	,
(	10888	)	,
(	10884	)	,
(	10880	)	,
(	10876	)	,
(	10872	)	,
(	10868	)	,
(	10864	)	,
(	10860	)	,
(	10856	)	,
(	10852	)	,
(	10848	)	,
(	10844	)	,
(	10840	)	,
(	10836	)	,
(	10832	)	,
(	10828	)	,
(	10824	)	,
(	10820	)	,
(	10816	)	,
(	10812	)	,
(	10808	)	,
(	10804	)	,
(	10800	)	,
(	10796	)	,
(	10792	)	,
(	10788	)	,
(	10784	)	,
(	10780	)	,
(	10776	)	,
(	10772	)	,
(	10768	)	,
(	10764	)	,
(	10760	)	,
(	10756	)	,
(	10752	)	,
(	10748	)	,
(	10744	)	,
(	10740	)	,
(	10736	)	,
(	10732	)	,
(	10728	)	,
(	10724	)	,
(	10720	)	,
(	10716	)	,
(	10712	)	,
(	10708	)	,
(	10704	)	,
(	10700	)	,
(	10696	)	,
(	10692	)	,
(	10688	)	,
(	10684	)	,
(	10680	)	,
(	10676	)	,
(	10672	)	,
(	10668	)	,
(	10664	)	,
(	10660	)	,
(	10656	)	,
(	10652	)	,
(	10648	)	,
(	10644	)	,
(	10640	)	,
(	10636	)	,
(	10632	)	,
(	10628	)	,
(	10624	)	,
(	10620	)	,
(	10616	)	,
(	10612	)	,
(	10608	)	,
(	10604	)	,
(	10600	)	,
(	10596	)	,
(	10592	)	,
(	10588	)	,
(	10584	)	,
(	10580	)	,
(	10576	)	,
(	10572	)	,
(	10568	)	,
(	10564	)	,
(	10560	)	,
(	10556	)	,
(	10552	)	,
(	10548	)	,
(	10544	)	,
(	10540	)	,
(	10536	)	,
(	10532	)	,
(	10528	)	,
(	10524	)	,
(	10520	)	,
(	10516	)	,
(	10512	)	,
(	10508	)	,
(	10504	)	,
(	10500	)	,
(	10496	)	,
(	10492	)	,
(	10488	)	,
(	10484	)	,
(	10480	)	,
(	10476	)	,
(	10472	)	,
(	10468	)	,
(	10464	)	,
(	10460	)	,
(	10456	)	,
(	10452	)	,
(	10448	)	,
(	10444	)	,
(	10440	)	,
(	10436	)	,
(	10432	)	,
(	10428	)	,
(	10424	)	,
(	10420	)	,
(	10416	)	,
(	10412	)	,
(	10408	)	,
(	10404	)	,
(	10400	)	,
(	10396	)	,
(	10392	)	,
(	10388	)	,
(	10384	)	,
(	10380	)	,
(	10376	)	,
(	10372	)	,
(	10368	)	,
(	10364	)	,
(	10360	)	,
(	10356	)	,
(	10352	)	,
(	10348	)	,
(	10344	)	,
(	10340	)	,
(	10336	)	,
(	10332	)	,
(	10328	)	,
(	10324	)	,
(	10320	)	,
(	10316	)	,
(	10312	)	,
(	10308	)	,
(	10304	)	,
(	10300	)	,
(	10296	)	,
(	10292	)	,
(	10288	)	,
(	10284	)	,
(	10280	)	,
(	10276	)	,
(	10272	)	,
(	10268	)	,
(	10264	)	,
(	10260	)	,
(	10256	)	,
(	10252	)	,
(	10248	)	,
(	10244	)	,
(	10240	)	,
(	10236	)	,
(	10232	)	,
(	10228	)	,
(	10224	)	,
(	10220	)	,
(	10216	)	,
(	10212	)	,
(	10208	)	,
(	10204	)	,
(	10200	)	,
(	10196	)	,
(	10192	)	,
(	10188	)	,
(	10184	)	,
(	10180	)	,
(	10176	)	,
(	10172	)	,
(	10168	)	,
(	10164	)	,
(	10160	)	,
(	10156	)	,
(	10152	)	,
(	10148	)	,
(	10144	)	,
(	10140	)	,
(	10136	)	,
(	10132	)	,
(	10128	)	,
(	10124	)	,
(	10120	)	,
(	10116	)	,
(	10112	)	,
(	10108	)	,
(	10104	)	,
(	10100	)	,
(	10096	)	,
(	10092	)	,
(	10088	)	,
(	10084	)	,
(	10080	)	,
(	10076	)	,
(	10072	)	,
(	10068	)	,
(	10064	)	,
(	10060	)	,
(	10056	)	,
(	10052	)	,
(	10048	)	,
(	10044	)	,
(	10040	)	,
(	10036	)	,
(	10032	)	,
(	10028	)	,
(	10024	)	,
(	10020	)	,
(	10016	)	,
(	10012	)	,
(	10008	)	,
(	10004	)	,
(	10000	)	,
(	9996	)	,
(	9992	)	,
(	9988	)	,
(	9984	)	,
(	9980	)	,
(	9976	)	,
(	9972	)	,
(	9968	)	,
(	9964	)	,
(	9960	)	,
(	9956	)	,
(	9952	)	,
(	9948	)	,
(	9944	)	,
(	9940	)	,
(	9936	)	,
(	9932	)	,
(	9928	)	,
(	9924	)	,
(	9920	)	,
(	9916	)	,
(	9912	)	,
(	9908	)	,
(	9904	)	,
(	9900	)	,
(	9896	)	,
(	9892	)	,
(	9888	)	,
(	9884	)	,
(	9880	)	,
(	9876	)	,
(	9872	)	,
(	9868	)	,
(	9864	)	,
(	9860	)	,
(	9856	)	,
(	9852	)	,
(	9848	)	,
(	9844	)	,
(	9840	)	,
(	9836	)	,
(	9832	)	,
(	9828	)	,
(	9824	)	,
(	9820	)	,
(	9816	)	,
(	9812	)	,
(	9808	)	,
(	9804	)	,
(	9800	)	,
(	9796	)	,
(	9792	)	,
(	9788	)	,
(	9784	)	,
(	9780	)	,
(	9776	)	,
(	9772	)	,
(	9768	)	,
(	9764	)	,
(	9760	)	,
(	9756	)	,
(	9752	)	,
(	9748	)	,
(	9744	)	,
(	9740	)	,
(	9736	)	,
(	9732	)	,
(	9728	)	,
(	9724	)	,
(	9720	)	,
(	9716	)	,
(	9712	)	,
(	9708	)	,
(	9704	)	,
(	9700	)	,
(	9696	)	,
(	9692	)	,
(	9688	)	,
(	9684	)	,
(	9680	)	,
(	9676	)	,
(	9672	)	,
(	9668	)	,
(	9664	)	,
(	9660	)	,
(	9656	)	,
(	9652	)	,
(	9648	)	,
(	9644	)	,
(	9640	)	,
(	9636	)	,
(	9632	)	,
(	9628	)	,
(	9624	)	,
(	9620	)	,
(	9616	)	,
(	9612	)	,
(	9608	)	,
(	9604	)	,
(	9600	)	,
(	9596	)	,
(	9592	)	,
(	9588	)	,
(	9584	)	,
(	9580	)	,
(	9576	)	,
(	9572	)	,
(	9568	)	,
(	9564	)	,
(	9560	)	,
(	9556	)	,
(	9552	)	,
(	9548	)	,
(	9544	)	,
(	9540	)	,
(	9536	)	,
(	9532	)	,
(	9528	)	,
(	9524	)	,
(	9520	)	,
(	9516	)	,
(	9512	)	,
(	9508	)	,
(	9504	)	,
(	9500	)	,
(	9496	)	,
(	9492	)	,
(	9488	)	,
(	9484	)	,
(	9480	)	,
(	9476	)	,
(	9472	)	,
(	9468	)	,
(	9464	)	,
(	9460	)	,
(	9456	)	,
(	9452	)	,
(	9448	)	,
(	9444	)	,
(	9440	)	,
(	9436	)	,
(	9432	)	,
(	9428	)	,
(	9424	)	,
(	9420	)	,
(	9416	)	,
(	9412	)	,
(	9408	)	,
(	9404	)	,
(	9400	)	,
(	9396	)	,
(	9392	)	,
(	9388	)	,
(	9384	)	,
(	9380	)	,
(	9376	)	,
(	9372	)	,
(	9368	)	,
(	9364	)	,
(	9360	)	,
(	9356	)	,
(	9352	)	,
(	9348	)	,
(	9344	)	,
(	9340	)	,
(	9336	)	,
(	9332	)	,
(	9328	)	,
(	9324	)	,
(	9320	)	,
(	9316	)	,
(	9312	)	,
(	9308	)	,
(	9304	)	,
(	9300	)	,
(	9296	)	,
(	9292	)	,
(	9288	)	,
(	9284	)	,
(	9280	)	,
(	9276	)	,
(	9272	)	,
(	9268	)	,
(	9264	)	,
(	9260	)	,
(	9256	)	,
(	9252	)	,
(	9248	)	,
(	9244	)	,
(	9240	)	,
(	9236	)	,
(	9232	)	,
(	9228	)	,
(	9224	)	,
(	9220	)	,
(	9216	)	,
(	9212	)	,
(	9208	)	,
(	9204	)	,
(	9200	)	,
(	9196	)	,
(	9192	)	,
(	9188	)	,
(	9184	)	,
(	9180	)	,
(	9176	)	,
(	9172	)	,
(	9168	)	,
(	9164	)	,
(	9160	)	,
(	9156	)	,
(	9152	)	,
(	9148	)	,
(	9144	)	,
(	9140	)	,
(	9136	)	,
(	9132	)	,
(	9128	)	,
(	9124	)	,
(	9120	)	,
(	9116	)	,
(	9112	)	,
(	9108	)	,
(	9104	)	,
(	9100	)	,
(	9096	)	,
(	9092	)	,
(	9088	)	,
(	9084	)	,
(	9080	)	,
(	9076	)	,
(	9072	)	,
(	9068	)	,
(	9064	)	,
(	9060	)	,
(	9056	)	,
(	9052	)	,
(	9048	)	,
(	9044	)	,
(	9040	)	,
(	9036	)	,
(	9032	)	,
(	9028	)	,
(	9024	)	,
(	9020	)	,
(	9016	)	,
(	9012	)	,
(	9008	)	,
(	9004	)	,
(	9000	)	,
(	8996	)	,
(	8992	)	,
(	8988	)	,
(	8984	)	,
(	8980	)	,
(	8976	)	,
(	8972	)	,
(	8968	)	,
(	8964	)	,
(	8960	)	,
(	8956	)	,
(	8952	)	,
(	8948	)	,
(	8944	)	,
(	8940	)	,
(	8936	)	,
(	8932	)	,
(	8928	)	,
(	8924	)	,
(	8920	)	,
(	8916	)	,
(	8912	)	,
(	8908	)	,
(	8904	)	,
(	8900	)	,
(	8896	)	,
(	8892	)	,
(	8888	)	,
(	8884	)	,
(	8880	)	,
(	8876	)	,
(	8872	)	,
(	8868	)	,
(	8864	)	,
(	8860	)	,
(	8856	)	,
(	8852	)	,
(	8848	)	,
(	8844	)	,
(	8840	)	,
(	8836	)	,
(	8832	)	,
(	8828	)	,
(	8824	)	,
(	8820	)	,
(	8816	)	,
(	8812	)	,
(	8808	)	,
(	8804	)	,
(	8800	)	,
(	8796	)	,
(	8792	)	,
(	8788	)	,
(	8784	)	,
(	8780	)	,
(	8776	)	,
(	8772	)	,
(	8768	)	,
(	8764	)	,
(	8760	)	,
(	8756	)	,
(	8752	)	,
(	8748	)	,
(	8744	)	,
(	8740	)	,
(	8736	)	,
(	8732	)	,
(	8728	)	,
(	8724	)	,
(	8720	)	,
(	8716	)	,
(	8712	)	,
(	8708	)	,
(	8704	)	,
(	8700	)	,
(	8696	)	,
(	8692	)	,
(	8688	)	,
(	8684	)	,
(	8680	)	,
(	8676	)	,
(	8672	)	,
(	8668	)	,
(	8664	)	,
(	8660	)	,
(	8656	)	,
(	8652	)	,
(	8648	)	,
(	8644	)	,
(	8640	)	,
(	8636	)	,
(	8632	)	,
(	8628	)	,
(	8624	)	,
(	8620	)	,
(	8616	)	,
(	8612	)	,
(	8608	)	,
(	8604	)	,
(	8600	)	,
(	8596	)	,
(	8592	)	,
(	8588	)	,
(	8584	)	,
(	8580	)	,
(	8576	)	,
(	8572	)	,
(	8568	)	,
(	8564	)	,
(	8560	)	,
(	8556	)	,
(	8552	)	,
(	8548	)	,
(	8544	)	,
(	8540	)	,
(	8536	)	,
(	8532	)	,
(	8528	)	,
(	8524	)	,
(	8520	)	,
(	8516	)	,
(	8512	)	,
(	8508	)	,
(	8504	)	,
(	8500	)	,
(	8496	)	,
(	8492	)	,
(	8488	)	,
(	8484	)	,
(	8480	)	,
(	8476	)	,
(	8472	)	,
(	8468	)	,
(	8464	)	,
(	8460	)	,
(	8456	)	,
(	8452	)	,
(	8448	)	,
(	8444	)	,
(	8440	)	,
(	8436	)	,
(	8432	)	,
(	8428	)	,
(	8424	)	,
(	8420	)	,
(	8416	)	,
(	8412	)	,
(	8408	)	,
(	8404	)	,
(	8400	)	,
(	8396	)	,
(	8392	)	,
(	8388	)	,
(	8384	)	,
(	8380	)	,
(	8376	)	,
(	8372	)	,
(	8368	)	,
(	8364	)	,
(	8360	)	,
(	8356	)	,
(	8352	)	,
(	8348	)	,
(	8344	)	,
(	8340	)	,
(	8336	)	,
(	8332	)	,
(	8328	)	,
(	8324	)	,
(	8320	)	,
(	8316	)	,
(	8312	)	,
(	8308	)	,
(	8304	)	,
(	8300	)	,
(	8296	)	,
(	8292	)	,
(	8288	)	,
(	8284	)	,
(	8280	)	,
(	8276	)	,
(	8272	)	,
(	8268	)	,
(	8264	)	,
(	8260	)	,
(	8256	)	,
(	8252	)	,
(	8248	)	,
(	8244	)	,
(	8240	)	,
(	8236	)	,
(	8232	)	,
(	8228	)	,
(	8224	)	,
(	8220	)	,
(	8216	)	,
(	8212	)	,
(	8208	)	,
(	8204	)	,
(	8200	)	,
(	8196	)	,
(	8192	)	,
(	8188	)	,
(	8184	)	,
(	8180	)	,
(	8176	)	,
(	8172	)	,
(	8168	)	,
(	8164	)	,
(	8160	)	,
(	8156	)	,
(	8152	)	,
(	8148	)	,
(	8144	)	,
(	8140	)	,
(	8136	)	,
(	8132	)	,
(	8128	)	,
(	8124	)	,
(	8120	)	,
(	8116	)	,
(	8112	)	,
(	8108	)	,
(	8104	)	,
(	8100	)	,
(	8096	)	,
(	8092	)	,
(	8088	)	,
(	8084	)	,
(	8080	)	,
(	8076	)	,
(	8072	)	,
(	8068	)	,
(	8064	)	,
(	8060	)	,
(	8056	)	,
(	8052	)	,
(	8048	)	,
(	8044	)	,
(	8040	)	,
(	8036	)	,
(	8032	)	,
(	8028	)	,
(	8024	)	,
(	8020	)	,
(	8016	)	,
(	8012	)	,
(	8008	)	,
(	8004	)	,
(	8000	)	,
(	7996	)	,
(	7992	)	,
(	7988	)	,
(	7984	)	,
(	7980	)	,
(	7976	)	,
(	7972	)	,
(	7968	)	,
(	7964	)	,
(	7960	)	,
(	7956	)	,
(	7952	)	,
(	7948	)	,
(	7944	)	,
(	7940	)	,
(	7936	)	,
(	7932	)	,
(	7928	)	,
(	7924	)	,
(	7920	)	,
(	7916	)	,
(	7912	)	,
(	7908	)	,
(	7904	)	,
(	7900	)	,
(	7896	)	,
(	7892	)	,
(	7888	)	,
(	7884	)	,
(	7880	)	,
(	7876	)	,
(	7872	)	,
(	7868	)	,
(	7864	)	,
(	7860	)	,
(	7856	)	,
(	7852	)	,
(	7848	)	,
(	7844	)	,
(	7840	)	,
(	7836	)	,
(	7832	)	,
(	7828	)	,
(	7824	)	,
(	7820	)	,
(	7816	)	,
(	7812	)	,
(	7808	)	,
(	7804	)	,
(	7800	)	,
(	7796	)	,
(	7792	)	,
(	7788	)	,
(	7784	)	,
(	7780	)	,
(	7776	)	,
(	7772	)	,
(	7768	)	,
(	7764	)	,
(	7760	)	,
(	7756	)	,
(	7752	)	,
(	7748	)	,
(	7744	)	,
(	7740	)	,
(	7736	)	,
(	7732	)	,
(	7728	)	,
(	7724	)	,
(	7720	)	,
(	7716	)	,
(	7712	)	,
(	7708	)	,
(	7704	)	,
(	7700	)	,
(	7696	)	,
(	7692	)	,
(	7688	)	,
(	7684	)	,
(	7680	)	,
(	7676	)	,
(	7672	)	,
(	7668	)	,
(	7664	)	,
(	7660	)	,
(	7656	)	,
(	7652	)	,
(	7648	)	,
(	7644	)	,
(	7640	)	,
(	7636	)	,
(	7632	)	,
(	7628	)	,
(	7624	)	,
(	7620	)	,
(	7616	)	,
(	7612	)	,
(	7608	)	,
(	7604	)	,
(	7600	)	,
(	7596	)	,
(	7592	)	,
(	7588	)	,
(	7584	)	,
(	7580	)	,
(	7576	)	,
(	7572	)	,
(	7568	)	,
(	7564	)	,
(	7560	)	,
(	7556	)	,
(	7552	)	,
(	7548	)	,
(	7544	)	,
(	7540	)	,
(	7536	)	,
(	7532	)	,
(	7528	)	,
(	7524	)	,
(	7520	)	,
(	7516	)	,
(	7512	)	,
(	7508	)	,
(	7504	)	,
(	7500	)	,
(	7496	)	,
(	7492	)	,
(	7488	)	,
(	7484	)	,
(	7480	)	,
(	7476	)	,
(	7472	)	,
(	7468	)	,
(	7464	)	,
(	7460	)	,
(	7456	)	,
(	7452	)	,
(	7448	)	,
(	7444	)	,
(	7440	)	,
(	7436	)	,
(	7432	)	,
(	7428	)	,
(	7424	)	,
(	7420	)	,
(	7416	)	,
(	7412	)	,
(	7408	)	,
(	7404	)	,
(	7400	)	,
(	7396	)	,
(	7392	)	,
(	7388	)	,
(	7384	)	,
(	7380	)	,
(	7376	)	,
(	7372	)	,
(	7368	)	,
(	7364	)	,
(	7360	)	,
(	7356	)	,
(	7352	)	,
(	7348	)	,
(	7344	)	,
(	7340	)	,
(	7336	)	,
(	7332	)	,
(	7328	)	,
(	7324	)	,
(	7320	)	,
(	7316	)	,
(	7312	)	,
(	7308	)	,
(	7304	)	,
(	7300	)	,
(	7296	)	,
(	7292	)	,
(	7288	)	,
(	7284	)	,
(	7280	)	,
(	7276	)	,
(	7272	)	,
(	7268	)	,
(	7264	)	,
(	7260	)	,
(	7256	)	,
(	7252	)	,
(	7248	)	,
(	7244	)	,
(	7240	)	,
(	7236	)	,
(	7232	)	,
(	7228	)	,
(	7224	)	,
(	7220	)	,
(	7216	)	,
(	7212	)	,
(	7208	)	,
(	7204	)	,
(	7200	)	,
(	7196	)	,
(	7192	)	,
(	7188	)	,
(	7184	)	,
(	7180	)	,
(	7176	)	,
(	7172	)	,
(	7168	)	,
(	7164	)	,
(	7160	)	,
(	7156	)	,
(	7152	)	,
(	7148	)	,
(	7144	)	,
(	7140	)	,
(	7136	)	,
(	7132	)	,
(	7128	)	,
(	7124	)	,
(	7120	)	,
(	7116	)	,
(	7112	)	,
(	7108	)	,
(	7104	)	,
(	7100	)	,
(	7096	)	,
(	7092	)	,
(	7088	)	,
(	7084	)	,
(	7080	)	,
(	7076	)	,
(	7072	)	,
(	7068	)	,
(	7064	)	,
(	7060	)	,
(	7056	)	,
(	7052	)	,
(	7048	)	,
(	7044	)	,
(	7040	)	,
(	7036	)	,
(	7032	)	,
(	7028	)	,
(	7024	)	,
(	7020	)	,
(	7016	)	,
(	7012	)	,
(	7008	)	,
(	7004	)	,
(	7000	)	,
(	6996	)	,
(	6992	)	,
(	6988	)	,
(	6984	)	,
(	6980	)	,
(	6976	)	,
(	6972	)	,
(	6968	)	,
(	6964	)	,
(	6960	)	,
(	6956	)	,
(	6952	)	,
(	6948	)	,
(	6944	)	,
(	6940	)	,
(	6936	)	,
(	6932	)	,
(	6928	)	,
(	6924	)	,
(	6920	)	,
(	6916	)	,
(	6912	)	,
(	6908	)	,
(	6904	)	,
(	6900	)	,
(	6896	)	,
(	6892	)	,
(	6888	)	,
(	6884	)	,
(	6880	)	,
(	6876	)	,
(	6872	)	,
(	6868	)	,
(	6864	)	,
(	6860	)	,
(	6856	)	,
(	6852	)	,
(	6848	)	,
(	6844	)	,
(	6840	)	,
(	6836	)	,
(	6832	)	,
(	6828	)	,
(	6824	)	,
(	6820	)	,
(	6816	)	,
(	6812	)	,
(	6808	)	,
(	6804	)	,
(	6800	)	,
(	6796	)	,
(	6792	)	,
(	6788	)	,
(	6784	)	,
(	6780	)	,
(	6776	)	,
(	6772	)	,
(	6768	)	,
(	6764	)	,
(	6760	)	,
(	6756	)	,
(	6752	)	,
(	6748	)	,
(	6744	)	,
(	6740	)	,
(	6736	)	,
(	6732	)	,
(	6728	)	,
(	6724	)	,
(	6720	)	,
(	6716	)	,
(	6712	)	,
(	6708	)	,
(	6704	)	,
(	6700	)	,
(	6696	)	,
(	6692	)	,
(	6688	)	,
(	6684	)	,
(	6680	)	,
(	6676	)	,
(	6672	)	,
(	6668	)	,
(	6664	)	,
(	6660	)	,
(	6656	)	,
(	6652	)	,
(	6648	)	,
(	6644	)	,
(	6640	)	,
(	6636	)	,
(	6632	)	,
(	6628	)	,
(	6624	)	,
(	6620	)	,
(	6616	)	,
(	6612	)	,
(	6608	)	,
(	6604	)	,
(	6600	)	,
(	6596	)	,
(	6592	)	,
(	6588	)	,
(	6584	)	,
(	6580	)	,
(	6576	)	,
(	6572	)	,
(	6568	)	,
(	6564	)	,
(	6560	)	,
(	6556	)	,
(	6552	)	,
(	6548	)	,
(	6544	)	,
(	6540	)	,
(	6536	)	,
(	6532	)	,
(	6528	)	,
(	6524	)	,
(	6520	)	,
(	6516	)	,
(	6512	)	,
(	6508	)	,
(	6504	)	,
(	6500	)	,
(	6496	)	,
(	6492	)	,
(	6488	)	,
(	6484	)	,
(	6480	)	,
(	6476	)	,
(	6472	)	,
(	6468	)	,
(	6464	)	,
(	6460	)	,
(	6456	)	,
(	6452	)	,
(	6448	)	,
(	6444	)	,
(	6440	)	,
(	6436	)	,
(	6432	)	,
(	6428	)	,
(	6424	)	,
(	6420	)	,
(	6416	)	,
(	6412	)	,
(	6408	)	,
(	6404	)	,
(	6400	)	,
(	6396	)	,
(	6392	)	,
(	6388	)	,
(	6384	)	,
(	6380	)	,
(	6376	)	,
(	6372	)	,
(	6368	)	,
(	6364	)	,
(	6360	)	,
(	6356	)	,
(	6352	)	,
(	6348	)	,
(	6344	)	,
(	6340	)	,
(	6336	)	,
(	6332	)	,
(	6328	)	,
(	6324	)	,
(	6320	)	,
(	6316	)	,
(	6312	)	,
(	6308	)	,
(	6304	)	,
(	6300	)	,
(	6296	)	,
(	6292	)	,
(	6288	)	,
(	6284	)	,
(	6280	)	,
(	6276	)	,
(	6272	)	,
(	6268	)	,
(	6264	)	,
(	6260	)	,
(	6256	)	,
(	6252	)	,
(	6248	)	,
(	6244	)	,
(	6240	)	,
(	6236	)	,
(	6232	)	,
(	6228	)	,
(	6224	)	,
(	6220	)	,
(	6216	)	,
(	6212	)	,
(	6208	)	,
(	6204	)	,
(	6200	)	,
(	6196	)	,
(	6192	)	,
(	6188	)	,
(	6184	)	,
(	6180	)	,
(	6176	)	,
(	6172	)	,
(	6168	)	,
(	6164	)	,
(	6160	)	,
(	6156	)	,
(	6152	)	,
(	6148	)	,
(	6144	)	,
(	6140	)	,
(	6136	)	,
(	6132	)	,
(	6128	)	,
(	6124	)	,
(	6120	)	,
(	6116	)	,
(	6112	)	,
(	6108	)	,
(	6104	)	,
(	6100	)	,
(	6096	)	,
(	6092	)	,
(	6088	)	,
(	6084	)	,
(	6080	)	,
(	6076	)	,
(	6072	)	,
(	6068	)	,
(	6064	)	,
(	6060	)	,
(	6056	)	,
(	6052	)	,
(	6048	)	,
(	6044	)	,
(	6040	)	,
(	6036	)	,
(	6032	)	,
(	6028	)	,
(	6024	)	,
(	6020	)	,
(	6016	)	,
(	6012	)	,
(	6008	)	,
(	6004	)	,
(	6000	)	,
(	5996	)	,
(	5992	)	,
(	5988	)	,
(	5984	)	,
(	5980	)	,
(	5976	)	,
(	5972	)	,
(	5968	)	,
(	5964	)	,
(	5960	)	,
(	5956	)	,
(	5952	)	,
(	5948	)	,
(	5944	)	,
(	5940	)	,
(	5936	)	,
(	5932	)	,
(	5928	)	,
(	5924	)	,
(	5920	)	,
(	5916	)	,
(	5912	)	,
(	5908	)	,
(	5904	)	,
(	5900	)	,
(	5896	)	,
(	5892	)	,
(	5888	)	,
(	5884	)	,
(	5880	)	,
(	5876	)	,
(	5872	)	,
(	5868	)	,
(	5864	)	,
(	5860	)	,
(	5856	)	,
(	5852	)	,
(	5848	)	,
(	5844	)	,
(	5840	)	,
(	5836	)	,
(	5832	)	,
(	5828	)	,
(	5824	)	,
(	5820	)	,
(	5816	)	,
(	5812	)	,
(	5808	)	,
(	5804	)	,
(	5800	)	,
(	5796	)	,
(	5792	)	,
(	5788	)	,
(	5784	)	,
(	5780	)	,
(	5776	)	,
(	5772	)	,
(	5768	)	,
(	5764	)	,
(	5760	)	,
(	5756	)	,
(	5752	)	,
(	5748	)	,
(	5744	)	,
(	5740	)	,
(	5736	)	,
(	5732	)	,
(	5728	)	,
(	5724	)	,
(	5720	)	,
(	5716	)	,
(	5712	)	,
(	5708	)	,
(	5704	)	,
(	5700	)	,
(	5696	)	,
(	5692	)	,
(	5688	)	,
(	5684	)	,
(	5680	)	,
(	5676	)	,
(	5672	)	,
(	5668	)	,
(	5664	)	,
(	5660	)	,
(	5656	)	,
(	5652	)	,
(	5648	)	,
(	5644	)	,
(	5640	)	,
(	5636	)	,
(	5632	)	,
(	5628	)	,
(	5624	)	,
(	5620	)	,
(	5616	)	,
(	5612	)	,
(	5608	)	,
(	5604	)	,
(	5600	)	,
(	5596	)	,
(	5592	)	,
(	5588	)	,
(	5584	)	,
(	5580	)	,
(	5576	)	,
(	5572	)	,
(	5568	)	,
(	5564	)	,
(	5560	)	,
(	5556	)	,
(	5552	)	,
(	5548	)	,
(	5544	)	,
(	5540	)	,
(	5536	)	,
(	5532	)	,
(	5528	)	,
(	5524	)	,
(	5520	)	,
(	5516	)	,
(	5512	)	,
(	5508	)	,
(	5504	)	,
(	5500	)	,
(	5496	)	,
(	5492	)	,
(	5488	)	,
(	5484	)	,
(	5480	)	,
(	5476	)	,
(	5472	)	,
(	5468	)	,
(	5464	)	,
(	5460	)	,
(	5456	)	,
(	5452	)	,
(	5448	)	,
(	5444	)	,
(	5440	)	,
(	5436	)	,
(	5432	)	,
(	5428	)	,
(	5424	)	,
(	5420	)	,
(	5416	)	,
(	5412	)	,
(	5408	)	,
(	5404	)	,
(	5400	)	,
(	5396	)	,
(	5392	)	,
(	5388	)	,
(	5384	)	,
(	5380	)	,
(	5376	)	,
(	5372	)	,
(	5368	)	,
(	5364	)	,
(	5360	)	,
(	5356	)	,
(	5352	)	,
(	5348	)	,
(	5344	)	,
(	5340	)	,
(	5336	)	,
(	5332	)	,
(	5328	)	,
(	5324	)	,
(	5320	)	,
(	5316	)	,
(	5312	)	,
(	5308	)	,
(	5304	)	,
(	5300	)	,
(	5296	)	,
(	5292	)	,
(	5288	)	,
(	5284	)	,
(	5280	)	,
(	5276	)	,
(	5272	)	,
(	5268	)	,
(	5264	)	,
(	5260	)	,
(	5256	)	,
(	5252	)	,
(	5248	)	,
(	5244	)	,
(	5240	)	,
(	5236	)	,
(	5232	)	,
(	5228	)	,
(	5224	)	,
(	5220	)	,
(	5216	)	,
(	5212	)	,
(	5208	)	,
(	5204	)	,
(	5200	)	,
(	5196	)	,
(	5192	)	,
(	5188	)	,
(	5184	)	,
(	5180	)	,
(	5176	)	,
(	5172	)	,
(	5168	)	,
(	5164	)	,
(	5160	)	,
(	5156	)	,
(	5152	)	,
(	5148	)	,
(	5144	)	,
(	5140	)	,
(	5136	)	,
(	5132	)	,
(	5128	)	,
(	5124	)	,
(	5120	)	,
(	5116	)	,
(	5112	)	,
(	5108	)	,
(	5104	)	,
(	5100	)	,
(	5096	)	,
(	5092	)	,
(	5088	)	,
(	5084	)	,
(	5080	)	,
(	5076	)	,
(	5072	)	,
(	5068	)	,
(	5064	)	,
(	5060	)	,
(	5056	)	,
(	5052	)	,
(	5048	)	,
(	5044	)	,
(	5040	)	,
(	5036	)	,
(	5032	)	,
(	5028	)	,
(	5024	)	,
(	5020	)	,
(	5016	)	,
(	5012	)	,
(	5008	)	,
(	5004	)	,
(	5000	)	,
(	4996	)	,
(	4992	)	,
(	4988	)	,
(	4984	)	,
(	4980	)	,
(	4976	)	,
(	4972	)	,
(	4968	)	,
(	4964	)	,
(	4960	)	,
(	4956	)	,
(	4952	)	,
(	4948	)	,
(	4944	)	,
(	4940	)	,
(	4936	)	,
(	4932	)	,
(	4928	)	,
(	4924	)	,
(	4920	)	,
(	4916	)	,
(	4912	)	,
(	4908	)	,
(	4904	)	,
(	4900	)	,
(	4896	)	,
(	4892	)	,
(	4888	)	,
(	4884	)	,
(	4880	)	,
(	4876	)	,
(	4872	)	,
(	4868	)	,
(	4864	)	,
(	4860	)	,
(	4856	)	,
(	4852	)	,
(	4848	)	,
(	4844	)	,
(	4840	)	,
(	4836	)	,
(	4832	)	,
(	4828	)	,
(	4824	)	,
(	4820	)	,
(	4816	)	,
(	4812	)	,
(	4808	)	,
(	4804	)	,
(	4800	)	,
(	4796	)	,
(	4792	)	,
(	4788	)	,
(	4784	)	,
(	4780	)	,
(	4776	)	,
(	4772	)	,
(	4768	)	,
(	4764	)	,
(	4760	)	,
(	4756	)	,
(	4752	)	,
(	4748	)	,
(	4744	)	,
(	4740	)	,
(	4736	)	,
(	4732	)	,
(	4728	)	,
(	4724	)	,
(	4720	)	,
(	4716	)	,
(	4712	)	,
(	4708	)	,
(	4704	)	,
(	4700	)	,
(	4696	)	,
(	4692	)	,
(	4688	)	,
(	4684	)	,
(	4680	)	,
(	4676	)	,
(	4672	)	,
(	4668	)	,
(	4664	)	,
(	4660	)	,
(	4656	)	,
(	4652	)	,
(	4648	)	,
(	4644	)	,
(	4640	)	,
(	4636	)	,
(	4632	)	,
(	4628	)	,
(	4624	)	,
(	4620	)	,
(	4616	)	,
(	4612	)	,
(	4608	)	,
(	4604	)	,
(	4600	)	,
(	4596	)	,
(	4592	)	,
(	4588	)	,
(	4584	)	,
(	4580	)	,
(	4576	)	,
(	4572	)	,
(	4568	)	,
(	4564	)	,
(	4560	)	,
(	4556	)	,
(	4552	)	,
(	4548	)	,
(	4544	)	,
(	4540	)	,
(	4536	)	,
(	4532	)	,
(	4528	)	,
(	4524	)	,
(	4520	)	,
(	4516	)	,
(	4512	)	,
(	4508	)	,
(	4504	)	,
(	4500	)	,
(	4496	)	,
(	4492	)	,
(	4488	)	,
(	4484	)	,
(	4480	)	,
(	4476	)	,
(	4472	)	,
(	4468	)	,
(	4464	)	,
(	4460	)	,
(	4456	)	,
(	4452	)	,
(	4448	)	,
(	4444	)	,
(	4440	)	,
(	4436	)	,
(	4432	)	,
(	4428	)	,
(	4424	)	,
(	4420	)	,
(	4416	)	,
(	4412	)	,
(	4408	)	,
(	4404	)	,
(	4400	)	,
(	4396	)	,
(	4392	)	,
(	4388	)	,
(	4384	)	,
(	4380	)	,
(	4376	)	,
(	4372	)	,
(	4368	)	,
(	4364	)	,
(	4360	)	,
(	4356	)	,
(	4352	)	,
(	4348	)	,
(	4344	)	,
(	4340	)	,
(	4336	)	,
(	4332	)	,
(	4328	)	,
(	4324	)	,
(	4320	)	,
(	4316	)	,
(	4312	)	,
(	4308	)	,
(	4304	)	,
(	4300	)	,
(	4296	)	,
(	4292	)	,
(	4288	)	,
(	4284	)	,
(	4280	)	,
(	4276	)	,
(	4272	)	,
(	4268	)	,
(	4264	)	,
(	4260	)	,
(	4256	)	,
(	4252	)	,
(	4248	)	,
(	4244	)	,
(	4240	)	,
(	4236	)	,
(	4232	)	,
(	4228	)	,
(	4224	)	,
(	4220	)	,
(	4216	)	,
(	4212	)	,
(	4208	)	,
(	4204	)	,
(	4200	)	,
(	4196	)	,
(	4192	)	,
(	4188	)	,
(	4184	)	,
(	4180	)	,
(	4176	)	,
(	4172	)	,
(	4168	)	,
(	4164	)	,
(	4160	)	,
(	4156	)	,
(	4152	)	,
(	4148	)	,
(	4144	)	,
(	4140	)	,
(	4136	)	,
(	4132	)	,
(	4128	)	,
(	4124	)	,
(	4120	)	,
(	4116	)	,
(	4112	)	,
(	4108	)	,
(	4104	)	,
(	4100	)	,
(	4096	)	,
(	4092	)	,
(	4088	)	,
(	4084	)	,
(	4080	)	,
(	4076	)	,
(	4072	)	,
(	4068	)	,
(	4064	)	,
(	4060	)	,
(	4056	)	,
(	4052	)	,
(	4048	)	,
(	4044	)	,
(	4040	)	,
(	4036	)	,
(	4032	)	,
(	4028	)	,
(	4024	)	,
(	4020	)	,
(	4016	)	,
(	4012	)	,
(	4008	)	,
(	4004	)	,
(	4000	)	,
(	3996	)	,
(	3992	)	,
(	3988	)	,
(	3984	)	,
(	3980	)	,
(	3976	)	,
(	3972	)	,
(	3968	)	,
(	3964	)	,
(	3960	)	,
(	3956	)	,
(	3952	)	,
(	3948	)	,
(	3944	)	,
(	3940	)	,
(	3936	)	,
(	3932	)	,
(	3928	)	,
(	3924	)	,
(	3920	)	,
(	3916	)	,
(	3912	)	,
(	3908	)	,
(	3904	)	,
(	3900	)	,
(	3896	)	,
(	3892	)	,
(	3888	)	,
(	3884	)	,
(	3880	)	,
(	3876	)	,
(	3872	)	,
(	3868	)	,
(	3864	)	,
(	3860	)	,
(	3856	)	,
(	3852	)	,
(	3848	)	,
(	3844	)	,
(	3840	)	,
(	3836	)	,
(	3832	)	,
(	3828	)	,
(	3824	)	,
(	3820	)	,
(	3816	)	,
(	3812	)	,
(	3808	)	,
(	3804	)	,
(	3800	)	,
(	3796	)	,
(	3792	)	,
(	3788	)	,
(	3784	)	,
(	3780	)	,
(	3776	)	,
(	3772	)	,
(	3768	)	,
(	3764	)	,
(	3760	)	,
(	3756	)	,
(	3752	)	,
(	3748	)	,
(	3744	)	,
(	3740	)	,
(	3736	)	,
(	3732	)	,
(	3728	)	,
(	3724	)	,
(	3720	)	,
(	3716	)	,
(	3712	)	,
(	3708	)	,
(	3704	)	,
(	3700	)	,
(	3696	)	,
(	3692	)	,
(	3688	)	,
(	3684	)	,
(	3680	)	,
(	3676	)	,
(	3672	)	,
(	3668	)	,
(	3664	)	,
(	3660	)	,
(	3656	)	,
(	3652	)	,
(	3648	)	,
(	3644	)	,
(	3640	)	,
(	3636	)	,
(	3632	)	,
(	3628	)	,
(	3624	)	,
(	3620	)	,
(	3616	)	,
(	3612	)	,
(	3608	)	,
(	3604	)	,
(	3600	)	,
(	3596	)	,
(	3592	)	,
(	3588	)	,
(	3584	)	,
(	3580	)	,
(	3576	)	,
(	3572	)	,
(	3568	)	,
(	3564	)	,
(	3560	)	,
(	3556	)	,
(	3552	)	,
(	3548	)	,
(	3544	)	,
(	3540	)	,
(	3536	)	,
(	3532	)	,
(	3528	)	,
(	3524	)	,
(	3520	)	,
(	3516	)	,
(	3512	)	,
(	3508	)	,
(	3504	)	,
(	3500	)	,
(	3496	)	,
(	3492	)	,
(	3488	)	,
(	3484	)	,
(	3480	)	,
(	3476	)	,
(	3472	)	,
(	3468	)	,
(	3464	)	,
(	3460	)	,
(	3456	)	,
(	3452	)	,
(	3448	)	,
(	3444	)	,
(	3440	)	,
(	3436	)	,
(	3432	)	,
(	3428	)	,
(	3424	)	,
(	3420	)	,
(	3416	)	,
(	3412	)	,
(	3408	)	,
(	3404	)	,
(	3400	)	,
(	3396	)	,
(	3392	)	,
(	3388	)	,
(	3384	)	,
(	3380	)	,
(	3376	)	,
(	3372	)	,
(	3368	)	,
(	3364	)	,
(	3360	)	,
(	3356	)	,
(	3352	)	,
(	3348	)	,
(	3344	)	,
(	3340	)	,
(	3336	)	,
(	3332	)	,
(	3328	)	,
(	3324	)	,
(	3320	)	,
(	3316	)	,
(	3312	)	,
(	3308	)	,
(	3304	)	,
(	3300	)	,
(	3296	)	,
(	3292	)	,
(	3288	)	,
(	3284	)	,
(	3280	)	,
(	3276	)	,
(	3272	)	,
(	3268	)	,
(	3264	)	,
(	3260	)	,
(	3256	)	,
(	3252	)	,
(	3248	)	,
(	3244	)	,
(	3240	)	,
(	3236	)	,
(	3232	)	,
(	3228	)	,
(	3224	)	,
(	3220	)	,
(	3216	)	,
(	3212	)	,
(	3208	)	,
(	3204	)	,
(	3200	)	,
(	3196	)	,
(	3192	)	,
(	3188	)	,
(	3184	)	,
(	3180	)	,
(	3176	)	,
(	3172	)	,
(	3168	)	,
(	3164	)	,
(	3160	)	,
(	3156	)	,
(	3152	)	,
(	3148	)	,
(	3144	)	,
(	3140	)	,
(	3136	)	,
(	3132	)	,
(	3128	)	,
(	3124	)	,
(	3120	)	,
(	3116	)	,
(	3112	)	,
(	3108	)	,
(	3104	)	,
(	3100	)	,
(	3096	)	,
(	3092	)	,
(	3088	)	,
(	3084	)	,
(	3080	)	,
(	3076	)	,
(	3072	)	,
(	3068	)	,
(	3064	)	,
(	3060	)	,
(	3056	)	,
(	3052	)	,
(	3048	)	,
(	3044	)	,
(	3040	)	,
(	3036	)	,
(	3032	)	,
(	3028	)	,
(	3024	)	,
(	3020	)	,
(	3016	)	,
(	3012	)	,
(	3008	)	,
(	3004	)	,
(	3000	)	,
(	2996	)	,
(	2992	)	,
(	2988	)	,
(	2984	)	,
(	2980	)	,
(	2976	)	,
(	2972	)	,
(	2968	)	,
(	2964	)	,
(	2960	)	,
(	2956	)	,
(	2952	)	,
(	2948	)	,
(	2944	)	,
(	2940	)	,
(	2936	)	,
(	2932	)	,
(	2928	)	,
(	2924	)	,
(	2920	)	,
(	2916	)	,
(	2912	)	,
(	2908	)	,
(	2904	)	,
(	2900	)	,
(	2896	)	,
(	2892	)	,
(	2888	)	,
(	2884	)	,
(	2880	)	,
(	2876	)	,
(	2872	)	,
(	2868	)	,
(	2864	)	,
(	2860	)	,
(	2856	)	,
(	2852	)	,
(	2848	)	,
(	2844	)	,
(	2840	)	,
(	2836	)	,
(	2832	)	,
(	2828	)	,
(	2824	)	,
(	2820	)	,
(	2816	)	,
(	2812	)	,
(	2808	)	,
(	2804	)	,
(	2800	)	,
(	2796	)	,
(	2792	)	,
(	2788	)	,
(	2784	)	,
(	2780	)	,
(	2776	)	,
(	2772	)	,
(	2768	)	,
(	2764	)	,
(	2760	)	,
(	2756	)	,
(	2752	)	,
(	2748	)	,
(	2744	)	,
(	2740	)	,
(	2736	)	,
(	2732	)	,
(	2728	)	,
(	2724	)	,
(	2720	)	,
(	2716	)	,
(	2712	)	,
(	2708	)	,
(	2704	)	,
(	2700	)	,
(	2696	)	,
(	2692	)	,
(	2688	)	,
(	2684	)	,
(	2680	)	,
(	2676	)	,
(	2672	)	,
(	2668	)	,
(	2664	)	,
(	2660	)	,
(	2656	)	,
(	2652	)	,
(	2648	)	,
(	2644	)	,
(	2640	)	,
(	2636	)	,
(	2632	)	,
(	2628	)	,
(	2624	)	,
(	2620	)	,
(	2616	)	,
(	2612	)	,
(	2608	)	,
(	2604	)	,
(	2600	)	,
(	2596	)	,
(	2592	)	,
(	2588	)	,
(	2584	)	,
(	2580	)	,
(	2576	)	,
(	2572	)	,
(	2568	)	,
(	2564	)	,
(	2560	)	,
(	2556	)	,
(	2552	)	,
(	2548	)	,
(	2544	)	,
(	2540	)	,
(	2536	)	,
(	2532	)	,
(	2528	)	,
(	2524	)	,
(	2520	)	,
(	2516	)	,
(	2512	)	,
(	2508	)	,
(	2504	)	,
(	2500	)	,
(	2496	)	,
(	2492	)	,
(	2488	)	,
(	2484	)	,
(	2480	)	,
(	2476	)	,
(	2472	)	,
(	2468	)	,
(	2464	)	,
(	2460	)	,
(	2456	)	,
(	2452	)	,
(	2448	)	,
(	2444	)	,
(	2440	)	,
(	2436	)	,
(	2432	)	,
(	2428	)	,
(	2424	)	,
(	2420	)	,
(	2416	)	,
(	2412	)	,
(	2408	)	,
(	2404	)	,
(	2400	)	,
(	2396	)	,
(	2392	)	,
(	2388	)	,
(	2384	)	,
(	2380	)	,
(	2376	)	,
(	2372	)	,
(	2368	)	,
(	2364	)	,
(	2360	)	,
(	2356	)	,
(	2352	)	,
(	2348	)	,
(	2344	)	,
(	2340	)	,
(	2336	)	,
(	2332	)	,
(	2328	)	,
(	2324	)	,
(	2320	)	,
(	2316	)	,
(	2312	)	,
(	2308	)	,
(	2304	)	,
(	2300	)	,
(	2296	)	,
(	2292	)	,
(	2288	)	,
(	2284	)	,
(	2280	)	,
(	2276	)	,
(	2272	)	,
(	2268	)	,
(	2264	)	,
(	2260	)	,
(	2256	)	,
(	2252	)	,
(	2248	)	,
(	2244	)	,
(	2240	)	,
(	2236	)	,
(	2232	)	,
(	2228	)	,
(	2224	)	,
(	2220	)	,
(	2216	)	,
(	2212	)	,
(	2208	)	,
(	2204	)	,
(	2200	)	,
(	2196	)	,
(	2192	)	,
(	2188	)	,
(	2184	)	,
(	2180	)	,
(	2176	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2100	)	,
(	2096	)	,
(	2092	)	,
(	2088	)	,
(	2084	)	,
(	2080	)	,
(	2076	)	,
(	2072	)	,
(	2068	)	,
(	2064	)	,
(	2060	)	,
(	2056	)	,
(	2052	)	,
(	2048	)	,
(	2044	)	,
(	2040	)	,
(	2036	)	,
(	2032	)	,
(	2028	)	,
(	2024	)	,
(	2020	)	,
(	2016	)	,
(	2012	)	,
(	2008	)	,
(	2004	)	,
(	2000	)	,
(	1996	)	,
(	1992	)	,
(	1988	)	,
(	1984	)	,
(	1980	)	,
(	1976	)	,
(	1972	)	,
(	1968	)	,
(	1964	)	,
(	1960	)	,
(	1956	)	,
(	1952	)	,
(	1948	)	,
(	1944	)	,
(	1940	)	,
(	1936	)	,
(	1932	)	,
(	1928	)	,
(	1924	)	,
(	1920	)	,
(	1916	)	,
(	1912	)	,
(	1908	)	,
(	1904	)	,
(	1900	)	,
(	1896	)	,
(	1892	)	,
(	1888	)	,
(	1884	)	,
(	1880	)	,
(	1876	)	,
(	1872	)	,
(	1868	)	,
(	1864	)	,
(	1860	)	,
(	1856	)	,
(	1852	)	,
(	1848	)	,
(	1844	)	,
(	1840	)	,
(	1836	)	,
(	1832	)	,
(	1828	)	,
(	1824	)	,
(	1820	)	,
(	1816	)	,
(	1812	)	,
(	1808	)	,
(	1804	)	,
(	1800	)	,
(	1796	)	,
(	1792	)	,
(	1788	)	,
(	1784	)	,
(	1780	)	,
(	1776	)	,
(	1772	)	,
(	1768	)	,
(	1764	)	,
(	1760	)	,
(	1756	)	,
(	1752	)	,
(	1748	)	,
(	1744	)	,
(	1740	)	,
(	1736	)	,
(	1732	)	,
(	1728	)	,
(	1724	)	,
(	1720	)	,
(	1716	)	,
(	1712	)	,
(	1708	)	,
(	1704	)	,
(	1700	)	,
(	1696	)	,
(	1692	)	,
(	1688	)	,
(	1684	)	,
(	1680	)	,
(	1676	)	,
(	1672	)	,
(	1668	)	,
(	1664	)	,
(	1660	)	,
(	1656	)	,
(	1652	)	,
(	1648	)	,
(	1644	)	,
(	1640	)	,
(	1636	)	,
(	1632	)	,
(	1628	)	,
(	1624	)	,
(	1620	)	,
(	1616	)	,
(	1612	)	,
(	1608	)	,
(	1604	)	,
(	1600	)	,
(	1596	)	,
(	1592	)	,
(	1588	)	,
(	1584	)	,
(	1580	)	,
(	1576	)	,
(	1572	)	,
(	1568	)	,
(	1564	)	,
(	1560	)	,
(	1556	)	,
(	1552	)	,
(	1548	)	,
(	1544	)	,
(	1540	)	,
(	1536	)	,
(	1532	)	,
(	1528	)	,
(	1524	)	,
(	1520	)	,
(	1516	)	,
(	1512	)	,
(	1508	)	,
(	1504	)	,
(	1500	)	,
(	1496	)	,
(	1492	)	,
(	1488	)	,
(	1484	)	,
(	1480	)	,
(	1476	)	,
(	1472	)	,
(	1468	)	,
(	1464	)	,
(	1460	)	,
(	1456	)	,
(	1452	)	,
(	1448	)	,
(	1444	)	,
(	1440	)	,
(	1436	)	,
(	1432	)	,
(	1428	)	,
(	1424	)	,
(	1420	)	,
(	1416	)	,
(	1412	)	,
(	1408	)	,
(	1404	)	,
(	1400	)	,
(	1396	)	,
(	1392	)	,
(	1388	)	,
(	1384	)	,
(	1380	)	,
(	1376	)	,
(	1372	)	,
(	1368	)	,
(	1364	)	,
(	1360	)	,
(	1356	)	,
(	1352	)	,
(	1348	)	,
(	1344	)	,
(	1340	)	,
(	1336	)	,
(	1332	)	,
(	1328	)	,
(	1324	)	,
(	1320	)	,
(	1316	)	,
(	1312	)	,
(	1308	)	,
(	1304	)	,
(	1300	)	,
(	1296	)	,
(	1292	)	,
(	1288	)	,
(	1284	)	,
(	1280	)	,
(	1276	)	,
(	1272	)	,
(	1268	)	,
(	1264	)	,
(	1260	)	,
(	1256	)	,
(	1252	)	,
(	1248	)	,
(	1244	)	,
(	1240	)	,
(	1236	)	,
(	1232	)	,
(	1228	)	,
(	1224	)	,
(	1220	)	,
(	1216	)	,
(	1212	)	,
(	1208	)	,
(	1204	)	,
(	1200	)	,
(	1196	)	,
(	1192	)	,
(	1188	)	,
(	1184	)	,
(	1180	)	,
(	1176	)	,
(	1172	)	,
(	1168	)	,
(	1164	)	,
(	1160	)	,
(	1156	)	,
(	1152	)	,
(	1148	)	,
(	1144	)	,
(	1140	)	,
(	1136	)	,
(	1132	)	,
(	1128	)	,
(	1124	)	,
(	1120	)	
	
 );
 
 end package buzzer_LUT_pkg;