library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package buzzer_LUT_pkg is
 
 type my_array is array (4095 downto 0) of integer;
 constant DtoBP_LUT : my_array := ( -- can this be the same name as the one used for the display?
 
(	16656	)	,
(	16653	)	,
(	16650	)	,
(	16647	)	,
(	16644	)	,
(	16641	)	,
(	16638	)	,
(	16635	)	,
(	16632	)	,
(	16629	)	,
(	16626	)	,
(	16623	)	,
(	16620	)	,
(	16617	)	,
(	16614	)	,
(	16611	)	,
(	16608	)	,
(	16605	)	,
(	16602	)	,
(	16599	)	,
(	16596	)	,
(	16593	)	,
(	16590	)	,
(	16587	)	,
(	16584	)	,
(	16581	)	,
(	16578	)	,
(	16575	)	,
(	16572	)	,
(	16569	)	,
(	16566	)	,
(	16563	)	,
(	16560	)	,
(	16557	)	,
(	16554	)	,
(	16551	)	,
(	16548	)	,
(	16545	)	,
(	16542	)	,
(	16539	)	,
(	16536	)	,
(	16533	)	,
(	16530	)	,
(	16527	)	,
(	16524	)	,
(	16521	)	,
(	16518	)	,
(	16515	)	,
(	16512	)	,
(	16509	)	,
(	16506	)	,
(	16503	)	,
(	16500	)	,
(	16497	)	,
(	16494	)	,
(	16491	)	,
(	16488	)	,
(	16485	)	,
(	16482	)	,
(	16479	)	,
(	16476	)	,
(	16473	)	,
(	16470	)	,
(	16467	)	,
(	16464	)	,
(	16461	)	,
(	16458	)	,
(	16455	)	,
(	16452	)	,
(	16449	)	,
(	16446	)	,
(	16443	)	,
(	16440	)	,
(	16437	)	,
(	16434	)	,
(	16431	)	,
(	16428	)	,
(	16425	)	,
(	16422	)	,
(	16419	)	,
(	16416	)	,
(	16413	)	,
(	16410	)	,
(	16407	)	,
(	16404	)	,
(	16401	)	,
(	16398	)	,
(	16395	)	,
(	16392	)	,
(	16389	)	,
(	16386	)	,
(	16383	)	,
(	16380	)	,
(	16377	)	,
(	16374	)	,
(	16371	)	,
(	16368	)	,
(	16365	)	,
(	16362	)	,
(	16359	)	,
(	16356	)	,
(	16353	)	,
(	16350	)	,
(	16347	)	,
(	16344	)	,
(	16341	)	,
(	16338	)	,
(	16335	)	,
(	16332	)	,
(	16329	)	,
(	16326	)	,
(	16323	)	,
(	16320	)	,
(	16317	)	,
(	16314	)	,
(	16311	)	,
(	16308	)	,
(	16305	)	,
(	16302	)	,
(	16299	)	,
(	16296	)	,
(	16293	)	,
(	16290	)	,
(	16287	)	,
(	16284	)	,
(	16281	)	,
(	16278	)	,
(	16275	)	,
(	16272	)	,
(	16269	)	,
(	16266	)	,
(	16263	)	,
(	16260	)	,
(	16257	)	,
(	16254	)	,
(	16251	)	,
(	16248	)	,
(	16245	)	,
(	16242	)	,
(	16239	)	,
(	16236	)	,
(	16233	)	,
(	16230	)	,
(	16227	)	,
(	16224	)	,
(	16221	)	,
(	16218	)	,
(	16215	)	,
(	16212	)	,
(	16209	)	,
(	16206	)	,
(	16203	)	,
(	16200	)	,
(	16197	)	,
(	16194	)	,
(	16191	)	,
(	16188	)	,
(	16185	)	,
(	16182	)	,
(	16179	)	,
(	16176	)	,
(	16173	)	,
(	16170	)	,
(	16167	)	,
(	16164	)	,
(	16161	)	,
(	16158	)	,
(	16155	)	,
(	16152	)	,
(	16149	)	,
(	16146	)	,
(	16143	)	,
(	16140	)	,
(	16137	)	,
(	16134	)	,
(	16131	)	,
(	16128	)	,
(	16125	)	,
(	16122	)	,
(	16119	)	,
(	16116	)	,
(	16113	)	,
(	16110	)	,
(	16107	)	,
(	16104	)	,
(	16101	)	,
(	16098	)	,
(	16095	)	,
(	16092	)	,
(	16089	)	,
(	16086	)	,
(	16083	)	,
(	16080	)	,
(	16077	)	,
(	16074	)	,
(	16071	)	,
(	16068	)	,
(	16065	)	,
(	16062	)	,
(	16059	)	,
(	16056	)	,
(	16053	)	,
(	16050	)	,
(	16047	)	,
(	16044	)	,
(	16041	)	,
(	16038	)	,
(	16035	)	,
(	16032	)	,
(	16029	)	,
(	16026	)	,
(	16023	)	,
(	16020	)	,
(	16017	)	,
(	16014	)	,
(	16011	)	,
(	16008	)	,
(	16005	)	,
(	16002	)	,
(	15999	)	,
(	15996	)	,
(	15993	)	,
(	15990	)	,
(	15987	)	,
(	15984	)	,
(	15981	)	,
(	15978	)	,
(	15975	)	,
(	15972	)	,
(	15969	)	,
(	15966	)	,
(	15963	)	,
(	15960	)	,
(	15957	)	,
(	15954	)	,
(	15951	)	,
(	15948	)	,
(	15945	)	,
(	15942	)	,
(	15939	)	,
(	15936	)	,
(	15933	)	,
(	15930	)	,
(	15927	)	,
(	15924	)	,
(	15921	)	,
(	15918	)	,
(	15915	)	,
(	15912	)	,
(	15909	)	,
(	15906	)	,
(	15903	)	,
(	15900	)	,
(	15897	)	,
(	15894	)	,
(	15891	)	,
(	15888	)	,
(	15885	)	,
(	15882	)	,
(	15879	)	,
(	15876	)	,
(	15873	)	,
(	15870	)	,
(	15867	)	,
(	15864	)	,
(	15861	)	,
(	15858	)	,
(	15855	)	,
(	15852	)	,
(	15849	)	,
(	15846	)	,
(	15843	)	,
(	15840	)	,
(	15837	)	,
(	15834	)	,
(	15831	)	,
(	15828	)	,
(	15825	)	,
(	15822	)	,
(	15819	)	,
(	15816	)	,
(	15813	)	,
(	15810	)	,
(	15807	)	,
(	15804	)	,
(	15801	)	,
(	15798	)	,
(	15795	)	,
(	15792	)	,
(	15789	)	,
(	15786	)	,
(	15783	)	,
(	15780	)	,
(	15777	)	,
(	15774	)	,
(	15771	)	,
(	15768	)	,
(	15765	)	,
(	15762	)	,
(	15759	)	,
(	15756	)	,
(	15753	)	,
(	15750	)	,
(	15747	)	,
(	15744	)	,
(	15741	)	,
(	15738	)	,
(	15735	)	,
(	15732	)	,
(	15729	)	,
(	15726	)	,
(	15723	)	,
(	15720	)	,
(	15717	)	,
(	15714	)	,
(	15711	)	,
(	15708	)	,
(	15705	)	,
(	15702	)	,
(	15699	)	,
(	15696	)	,
(	15693	)	,
(	15690	)	,
(	15687	)	,
(	15684	)	,
(	15681	)	,
(	15678	)	,
(	15675	)	,
(	15672	)	,
(	15669	)	,
(	15666	)	,
(	15663	)	,
(	15660	)	,
(	15657	)	,
(	15654	)	,
(	15651	)	,
(	15648	)	,
(	15645	)	,
(	15642	)	,
(	15639	)	,
(	15636	)	,
(	15633	)	,
(	15630	)	,
(	15627	)	,
(	15624	)	,
(	15621	)	,
(	15618	)	,
(	15615	)	,
(	15612	)	,
(	15609	)	,
(	15606	)	,
(	15603	)	,
(	15600	)	,
(	15597	)	,
(	15594	)	,
(	15591	)	,
(	15588	)	,
(	15585	)	,
(	15582	)	,
(	15579	)	,
(	15576	)	,
(	15573	)	,
(	15570	)	,
(	15567	)	,
(	15564	)	,
(	15561	)	,
(	15558	)	,
(	15555	)	,
(	15552	)	,
(	15549	)	,
(	15546	)	,
(	15543	)	,
(	15540	)	,
(	15537	)	,
(	15534	)	,
(	15531	)	,
(	15528	)	,
(	15525	)	,
(	15522	)	,
(	15519	)	,
(	15516	)	,
(	15513	)	,
(	15510	)	,
(	15507	)	,
(	15504	)	,
(	15501	)	,
(	15498	)	,
(	15495	)	,
(	15492	)	,
(	15489	)	,
(	15486	)	,
(	15483	)	,
(	15480	)	,
(	15477	)	,
(	15474	)	,
(	15471	)	,
(	15468	)	,
(	15465	)	,
(	15462	)	,
(	15459	)	,
(	15456	)	,
(	15453	)	,
(	15450	)	,
(	15447	)	,
(	15444	)	,
(	15441	)	,
(	15438	)	,
(	15435	)	,
(	15432	)	,
(	15429	)	,
(	15426	)	,
(	15423	)	,
(	15420	)	,
(	15417	)	,
(	15414	)	,
(	15411	)	,
(	15408	)	,
(	15405	)	,
(	15402	)	,
(	15399	)	,
(	15396	)	,
(	15393	)	,
(	15390	)	,
(	15387	)	,
(	15384	)	,
(	15381	)	,
(	15378	)	,
(	15375	)	,
(	15372	)	,
(	15369	)	,
(	15366	)	,
(	15363	)	,
(	15360	)	,
(	15357	)	,
(	15354	)	,
(	15351	)	,
(	15348	)	,
(	15345	)	,
(	15342	)	,
(	15339	)	,
(	15336	)	,
(	15333	)	,
(	15330	)	,
(	15327	)	,
(	15324	)	,
(	15321	)	,
(	15318	)	,
(	15315	)	,
(	15312	)	,
(	15309	)	,
(	15306	)	,
(	15303	)	,
(	15300	)	,
(	15297	)	,
(	15294	)	,
(	15291	)	,
(	15288	)	,
(	15285	)	,
(	15282	)	,
(	15279	)	,
(	15276	)	,
(	15273	)	,
(	15270	)	,
(	15267	)	,
(	15264	)	,
(	15261	)	,
(	15258	)	,
(	15255	)	,
(	15252	)	,
(	15249	)	,
(	15246	)	,
(	15243	)	,
(	15240	)	,
(	15237	)	,
(	15234	)	,
(	15231	)	,
(	15228	)	,
(	15225	)	,
(	15222	)	,
(	15219	)	,
(	15216	)	,
(	15213	)	,
(	15210	)	,
(	15207	)	,
(	15204	)	,
(	15201	)	,
(	15198	)	,
(	15195	)	,
(	15192	)	,
(	15189	)	,
(	15186	)	,
(	15183	)	,
(	15180	)	,
(	15177	)	,
(	15174	)	,
(	15171	)	,
(	15168	)	,
(	15165	)	,
(	15162	)	,
(	15159	)	,
(	15156	)	,
(	15153	)	,
(	15150	)	,
(	15147	)	,
(	15144	)	,
(	15141	)	,
(	15138	)	,
(	15135	)	,
(	15132	)	,
(	15129	)	,
(	15126	)	,
(	15123	)	,
(	15120	)	,
(	15117	)	,
(	15114	)	,
(	15111	)	,
(	15108	)	,
(	15105	)	,
(	15102	)	,
(	15099	)	,
(	15096	)	,
(	15093	)	,
(	15090	)	,
(	15087	)	,
(	15084	)	,
(	15081	)	,
(	15078	)	,
(	15075	)	,
(	15072	)	,
(	15069	)	,
(	15066	)	,
(	15063	)	,
(	15060	)	,
(	15057	)	,
(	15054	)	,
(	15051	)	,
(	15048	)	,
(	15045	)	,
(	15042	)	,
(	15039	)	,
(	15036	)	,
(	15033	)	,
(	15030	)	,
(	15027	)	,
(	15024	)	,
(	15021	)	,
(	15018	)	,
(	15015	)	,
(	15012	)	,
(	15009	)	,
(	15006	)	,
(	15003	)	,
(	15000	)	,
(	14997	)	,
(	14994	)	,
(	14991	)	,
(	14988	)	,
(	14985	)	,
(	14982	)	,
(	14979	)	,
(	14976	)	,
(	14973	)	,
(	14970	)	,
(	14967	)	,
(	14964	)	,
(	14961	)	,
(	14958	)	,
(	14955	)	,
(	14952	)	,
(	14949	)	,
(	14946	)	,
(	14943	)	,
(	14940	)	,
(	14937	)	,
(	14934	)	,
(	14931	)	,
(	14928	)	,
(	14925	)	,
(	14922	)	,
(	14919	)	,
(	14916	)	,
(	14913	)	,
(	14910	)	,
(	14907	)	,
(	14904	)	,
(	14901	)	,
(	14898	)	,
(	14895	)	,
(	14892	)	,
(	14889	)	,
(	14886	)	,
(	14883	)	,
(	14880	)	,
(	14877	)	,
(	14874	)	,
(	14871	)	,
(	14868	)	,
(	14865	)	,
(	14862	)	,
(	14859	)	,
(	14856	)	,
(	14853	)	,
(	14850	)	,
(	14847	)	,
(	14844	)	,
(	14841	)	,
(	14838	)	,
(	14835	)	,
(	14832	)	,
(	14829	)	,
(	14826	)	,
(	14823	)	,
(	14820	)	,
(	14817	)	,
(	14814	)	,
(	14811	)	,
(	14808	)	,
(	14805	)	,
(	14802	)	,
(	14799	)	,
(	14796	)	,
(	14793	)	,
(	14790	)	,
(	14787	)	,
(	14784	)	,
(	14781	)	,
(	14778	)	,
(	14775	)	,
(	14772	)	,
(	14769	)	,
(	14766	)	,
(	14763	)	,
(	14760	)	,
(	14757	)	,
(	14754	)	,
(	14751	)	,
(	14748	)	,
(	14745	)	,
(	14742	)	,
(	14739	)	,
(	14736	)	,
(	14733	)	,
(	14730	)	,
(	14727	)	,
(	14724	)	,
(	14721	)	,
(	14718	)	,
(	14715	)	,
(	14712	)	,
(	14709	)	,
(	14706	)	,
(	14703	)	,
(	14700	)	,
(	14697	)	,
(	14694	)	,
(	14691	)	,
(	14688	)	,
(	14685	)	,
(	14682	)	,
(	14679	)	,
(	14676	)	,
(	14673	)	,
(	14670	)	,
(	14667	)	,
(	14664	)	,
(	14661	)	,
(	14658	)	,
(	14655	)	,
(	14652	)	,
(	14649	)	,
(	14646	)	,
(	14643	)	,
(	14640	)	,
(	14637	)	,
(	14634	)	,
(	14631	)	,
(	14628	)	,
(	14625	)	,
(	14622	)	,
(	14619	)	,
(	14616	)	,
(	14613	)	,
(	14610	)	,
(	14607	)	,
(	14604	)	,
(	14601	)	,
(	14598	)	,
(	14595	)	,
(	14592	)	,
(	14589	)	,
(	14586	)	,
(	14583	)	,
(	14580	)	,
(	14577	)	,
(	14574	)	,
(	14571	)	,
(	14568	)	,
(	14565	)	,
(	14562	)	,
(	14559	)	,
(	14556	)	,
(	14553	)	,
(	14550	)	,
(	14547	)	,
(	14544	)	,
(	14541	)	,
(	14538	)	,
(	14535	)	,
(	14532	)	,
(	14529	)	,
(	14526	)	,
(	14523	)	,
(	14520	)	,
(	14517	)	,
(	14514	)	,
(	14511	)	,
(	14508	)	,
(	14505	)	,
(	14502	)	,
(	14499	)	,
(	14496	)	,
(	14493	)	,
(	14490	)	,
(	14487	)	,
(	14484	)	,
(	14481	)	,
(	14478	)	,
(	14475	)	,
(	14472	)	,
(	14469	)	,
(	14466	)	,
(	14463	)	,
(	14460	)	,
(	14457	)	,
(	14454	)	,
(	14451	)	,
(	14448	)	,
(	14445	)	,
(	14442	)	,
(	14439	)	,
(	14436	)	,
(	14433	)	,
(	14430	)	,
(	14427	)	,
(	14424	)	,
(	14421	)	,
(	14418	)	,
(	14415	)	,
(	14412	)	,
(	14409	)	,
(	14406	)	,
(	14403	)	,
(	14400	)	,
(	14397	)	,
(	14394	)	,
(	14391	)	,
(	14388	)	,
(	14385	)	,
(	14382	)	,
(	14379	)	,
(	14376	)	,
(	14373	)	,
(	14370	)	,
(	14367	)	,
(	14364	)	,
(	14361	)	,
(	14358	)	,
(	14355	)	,
(	14352	)	,
(	14349	)	,
(	14346	)	,
(	14343	)	,
(	14340	)	,
(	14337	)	,
(	14334	)	,
(	14331	)	,
(	14328	)	,
(	14325	)	,
(	14322	)	,
(	14319	)	,
(	14316	)	,
(	14313	)	,
(	14310	)	,
(	14307	)	,
(	14304	)	,
(	14301	)	,
(	14298	)	,
(	14295	)	,
(	14292	)	,
(	14289	)	,
(	14286	)	,
(	14283	)	,
(	14280	)	,
(	14277	)	,
(	14274	)	,
(	14271	)	,
(	14268	)	,
(	14265	)	,
(	14262	)	,
(	14259	)	,
(	14256	)	,
(	14253	)	,
(	14250	)	,
(	14247	)	,
(	14244	)	,
(	14241	)	,
(	14238	)	,
(	14235	)	,
(	14232	)	,
(	14229	)	,
(	14226	)	,
(	14223	)	,
(	14220	)	,
(	14217	)	,
(	14214	)	,
(	14211	)	,
(	14208	)	,
(	14205	)	,
(	14202	)	,
(	14199	)	,
(	14196	)	,
(	14193	)	,
(	14190	)	,
(	14187	)	,
(	14184	)	,
(	14181	)	,
(	14178	)	,
(	14175	)	,
(	14172	)	,
(	14169	)	,
(	14166	)	,
(	14163	)	,
(	14160	)	,
(	14157	)	,
(	14154	)	,
(	14151	)	,
(	14148	)	,
(	14145	)	,
(	14142	)	,
(	14139	)	,
(	14136	)	,
(	14133	)	,
(	14130	)	,
(	14127	)	,
(	14124	)	,
(	14121	)	,
(	14118	)	,
(	14115	)	,
(	14112	)	,
(	14109	)	,
(	14106	)	,
(	14103	)	,
(	14100	)	,
(	14097	)	,
(	14094	)	,
(	14091	)	,
(	14088	)	,
(	14085	)	,
(	14082	)	,
(	14079	)	,
(	14076	)	,
(	14073	)	,
(	14070	)	,
(	14067	)	,
(	14064	)	,
(	14061	)	,
(	14058	)	,
(	14055	)	,
(	14052	)	,
(	14049	)	,
(	14046	)	,
(	14043	)	,
(	14040	)	,
(	14037	)	,
(	14034	)	,
(	14031	)	,
(	14028	)	,
(	14025	)	,
(	14022	)	,
(	14019	)	,
(	14016	)	,
(	14013	)	,
(	14010	)	,
(	14007	)	,
(	14004	)	,
(	14001	)	,
(	13998	)	,
(	13995	)	,
(	13992	)	,
(	13989	)	,
(	13986	)	,
(	13983	)	,
(	13980	)	,
(	13977	)	,
(	13974	)	,
(	13971	)	,
(	13968	)	,
(	13965	)	,
(	13962	)	,
(	13959	)	,
(	13956	)	,
(	13953	)	,
(	13950	)	,
(	13947	)	,
(	13944	)	,
(	13941	)	,
(	13938	)	,
(	13935	)	,
(	13932	)	,
(	13929	)	,
(	13926	)	,
(	13923	)	,
(	13920	)	,
(	13917	)	,
(	13914	)	,
(	13911	)	,
(	13908	)	,
(	13905	)	,
(	13902	)	,
(	13899	)	,
(	13896	)	,
(	13893	)	,
(	13890	)	,
(	13887	)	,
(	13884	)	,
(	13881	)	,
(	13878	)	,
(	13875	)	,
(	13872	)	,
(	13869	)	,
(	13866	)	,
(	13863	)	,
(	13860	)	,
(	13857	)	,
(	13854	)	,
(	13851	)	,
(	13848	)	,
(	13845	)	,
(	13842	)	,
(	13839	)	,
(	13836	)	,
(	13833	)	,
(	13830	)	,
(	13827	)	,
(	13824	)	,
(	13821	)	,
(	13818	)	,
(	13815	)	,
(	13812	)	,
(	13809	)	,
(	13806	)	,
(	13803	)	,
(	13800	)	,
(	13797	)	,
(	13794	)	,
(	13791	)	,
(	13788	)	,
(	13785	)	,
(	13782	)	,
(	13779	)	,
(	13776	)	,
(	13773	)	,
(	13770	)	,
(	13767	)	,
(	13764	)	,
(	13761	)	,
(	13758	)	,
(	13755	)	,
(	13752	)	,
(	13749	)	,
(	13746	)	,
(	13743	)	,
(	13740	)	,
(	13737	)	,
(	13734	)	,
(	13731	)	,
(	13728	)	,
(	13725	)	,
(	13722	)	,
(	13719	)	,
(	13716	)	,
(	13713	)	,
(	13710	)	,
(	13707	)	,
(	13704	)	,
(	13701	)	,
(	13698	)	,
(	13695	)	,
(	13692	)	,
(	13689	)	,
(	13686	)	,
(	13683	)	,
(	13680	)	,
(	13677	)	,
(	13674	)	,
(	13671	)	,
(	13668	)	,
(	13665	)	,
(	13662	)	,
(	13659	)	,
(	13656	)	,
(	13653	)	,
(	13650	)	,
(	13647	)	,
(	13644	)	,
(	13641	)	,
(	13638	)	,
(	13635	)	,
(	13632	)	,
(	13629	)	,
(	13626	)	,
(	13623	)	,
(	13620	)	,
(	13617	)	,
(	13614	)	,
(	13611	)	,
(	13608	)	,
(	13605	)	,
(	13602	)	,
(	13599	)	,
(	13596	)	,
(	13593	)	,
(	13590	)	,
(	13587	)	,
(	13584	)	,
(	13581	)	,
(	13578	)	,
(	13575	)	,
(	13572	)	,
(	13569	)	,
(	13566	)	,
(	13563	)	,
(	13560	)	,
(	13557	)	,
(	13554	)	,
(	13551	)	,
(	13548	)	,
(	13545	)	,
(	13542	)	,
(	13539	)	,
(	13536	)	,
(	13533	)	,
(	13530	)	,
(	13527	)	,
(	13524	)	,
(	13521	)	,
(	13518	)	,
(	13515	)	,
(	13512	)	,
(	13509	)	,
(	13506	)	,
(	13503	)	,
(	13500	)	,
(	13497	)	,
(	13494	)	,
(	13491	)	,
(	13488	)	,
(	13485	)	,
(	13482	)	,
(	13479	)	,
(	13476	)	,
(	13473	)	,
(	13470	)	,
(	13467	)	,
(	13464	)	,
(	13461	)	,
(	13458	)	,
(	13455	)	,
(	13452	)	,
(	13449	)	,
(	13446	)	,
(	13443	)	,
(	13440	)	,
(	13437	)	,
(	13434	)	,
(	13431	)	,
(	13428	)	,
(	13425	)	,
(	13422	)	,
(	13419	)	,
(	13416	)	,
(	13413	)	,
(	13410	)	,
(	13407	)	,
(	13404	)	,
(	13401	)	,
(	13398	)	,
(	13395	)	,
(	13392	)	,
(	13389	)	,
(	13386	)	,
(	13383	)	,
(	13380	)	,
(	13377	)	,
(	13374	)	,
(	13371	)	,
(	13368	)	,
(	13365	)	,
(	13362	)	,
(	13359	)	,
(	13356	)	,
(	13353	)	,
(	13350	)	,
(	13347	)	,
(	13344	)	,
(	13341	)	,
(	13338	)	,
(	13335	)	,
(	13332	)	,
(	13329	)	,
(	13326	)	,
(	13323	)	,
(	13320	)	,
(	13317	)	,
(	13314	)	,
(	13311	)	,
(	13308	)	,
(	13305	)	,
(	13302	)	,
(	13299	)	,
(	13296	)	,
(	13293	)	,
(	13290	)	,
(	13287	)	,
(	13284	)	,
(	13281	)	,
(	13278	)	,
(	13275	)	,
(	13272	)	,
(	13269	)	,
(	13266	)	,
(	13263	)	,
(	13260	)	,
(	13257	)	,
(	13254	)	,
(	13251	)	,
(	13248	)	,
(	13245	)	,
(	13242	)	,
(	13239	)	,
(	13236	)	,
(	13233	)	,
(	13230	)	,
(	13227	)	,
(	13224	)	,
(	13221	)	,
(	13218	)	,
(	13215	)	,
(	13212	)	,
(	13209	)	,
(	13206	)	,
(	13203	)	,
(	13200	)	,
(	13197	)	,
(	13194	)	,
(	13191	)	,
(	13188	)	,
(	13185	)	,
(	13182	)	,
(	13179	)	,
(	13176	)	,
(	13173	)	,
(	13170	)	,
(	13167	)	,
(	13164	)	,
(	13161	)	,
(	13158	)	,
(	13155	)	,
(	13152	)	,
(	13149	)	,
(	13146	)	,
(	13143	)	,
(	13140	)	,
(	13137	)	,
(	13134	)	,
(	13131	)	,
(	13128	)	,
(	13125	)	,
(	13122	)	,
(	13119	)	,
(	13116	)	,
(	13113	)	,
(	13110	)	,
(	13107	)	,
(	13104	)	,
(	13101	)	,
(	13098	)	,
(	13095	)	,
(	13092	)	,
(	13089	)	,
(	13086	)	,
(	13083	)	,
(	13080	)	,
(	13077	)	,
(	13074	)	,
(	13071	)	,
(	13068	)	,
(	13065	)	,
(	13062	)	,
(	13059	)	,
(	13056	)	,
(	13053	)	,
(	13050	)	,
(	13047	)	,
(	13044	)	,
(	13041	)	,
(	13038	)	,
(	13035	)	,
(	13032	)	,
(	13029	)	,
(	13026	)	,
(	13023	)	,
(	13020	)	,
(	13017	)	,
(	13014	)	,
(	13011	)	,
(	13008	)	,
(	13005	)	,
(	13002	)	,
(	12999	)	,
(	12996	)	,
(	12993	)	,
(	12990	)	,
(	12987	)	,
(	12984	)	,
(	12981	)	,
(	12978	)	,
(	12975	)	,
(	12972	)	,
(	12969	)	,
(	12966	)	,
(	12963	)	,
(	12960	)	,
(	12957	)	,
(	12954	)	,
(	12951	)	,
(	12948	)	,
(	12945	)	,
(	12942	)	,
(	12939	)	,
(	12936	)	,
(	12933	)	,
(	12930	)	,
(	12927	)	,
(	12924	)	,
(	12921	)	,
(	12918	)	,
(	12915	)	,
(	12912	)	,
(	12909	)	,
(	12906	)	,
(	12903	)	,
(	12900	)	,
(	12897	)	,
(	12894	)	,
(	12891	)	,
(	12888	)	,
(	12885	)	,
(	12882	)	,
(	12879	)	,
(	12876	)	,
(	12873	)	,
(	12870	)	,
(	12867	)	,
(	12864	)	,
(	12861	)	,
(	12858	)	,
(	12855	)	,
(	12852	)	,
(	12849	)	,
(	12846	)	,
(	12843	)	,
(	12840	)	,
(	12837	)	,
(	12834	)	,
(	12831	)	,
(	12828	)	,
(	12825	)	,
(	12822	)	,
(	12819	)	,
(	12816	)	,
(	12813	)	,
(	12810	)	,
(	12807	)	,
(	12804	)	,
(	12801	)	,
(	12798	)	,
(	12795	)	,
(	12792	)	,
(	12789	)	,
(	12786	)	,
(	12783	)	,
(	12780	)	,
(	12777	)	,
(	12774	)	,
(	12771	)	,
(	12768	)	,
(	12765	)	,
(	12762	)	,
(	12759	)	,
(	12756	)	,
(	12753	)	,
(	12750	)	,
(	12747	)	,
(	12744	)	,
(	12741	)	,
(	12738	)	,
(	12735	)	,
(	12732	)	,
(	12729	)	,
(	12726	)	,
(	12723	)	,
(	12720	)	,
(	12717	)	,
(	12714	)	,
(	12711	)	,
(	12708	)	,
(	12705	)	,
(	12702	)	,
(	12699	)	,
(	12696	)	,
(	12693	)	,
(	12690	)	,
(	12687	)	,
(	12684	)	,
(	12681	)	,
(	12678	)	,
(	12675	)	,
(	12672	)	,
(	12669	)	,
(	12666	)	,
(	12663	)	,
(	12660	)	,
(	12657	)	,
(	12654	)	,
(	12651	)	,
(	12648	)	,
(	12645	)	,
(	12642	)	,
(	12639	)	,
(	12636	)	,
(	12633	)	,
(	12630	)	,
(	12627	)	,
(	12624	)	,
(	12621	)	,
(	12618	)	,
(	12615	)	,
(	12612	)	,
(	12609	)	,
(	12606	)	,
(	12603	)	,
(	12600	)	,
(	12597	)	,
(	12594	)	,
(	12591	)	,
(	12588	)	,
(	12585	)	,
(	12582	)	,
(	12579	)	,
(	12576	)	,
(	12573	)	,
(	12570	)	,
(	12567	)	,
(	12564	)	,
(	12561	)	,
(	12558	)	,
(	12555	)	,
(	12552	)	,
(	12549	)	,
(	12546	)	,
(	12543	)	,
(	12540	)	,
(	12537	)	,
(	12534	)	,
(	12531	)	,
(	12528	)	,
(	12525	)	,
(	12522	)	,
(	12519	)	,
(	12516	)	,
(	12513	)	,
(	12510	)	,
(	12507	)	,
(	12504	)	,
(	12501	)	,
(	12498	)	,
(	12495	)	,
(	12492	)	,
(	12489	)	,
(	12486	)	,
(	12483	)	,
(	12480	)	,
(	12477	)	,
(	12474	)	,
(	12471	)	,
(	12468	)	,
(	12465	)	,
(	12462	)	,
(	12459	)	,
(	12456	)	,
(	12453	)	,
(	12450	)	,
(	12447	)	,
(	12444	)	,
(	12441	)	,
(	12438	)	,
(	12435	)	,
(	12432	)	,
(	12429	)	,
(	12426	)	,
(	12423	)	,
(	12420	)	,
(	12417	)	,
(	12414	)	,
(	12411	)	,
(	12408	)	,
(	12405	)	,
(	12402	)	,
(	12399	)	,
(	12396	)	,
(	12393	)	,
(	12390	)	,
(	12387	)	,
(	12384	)	,
(	12381	)	,
(	12378	)	,
(	12375	)	,
(	12372	)	,
(	12369	)	,
(	12366	)	,
(	12363	)	,
(	12360	)	,
(	12357	)	,
(	12354	)	,
(	12351	)	,
(	12348	)	,
(	12345	)	,
(	12342	)	,
(	12339	)	,
(	12336	)	,
(	12333	)	,
(	12330	)	,
(	12327	)	,
(	12324	)	,
(	12321	)	,
(	12318	)	,
(	12315	)	,
(	12312	)	,
(	12309	)	,
(	12306	)	,
(	12303	)	,
(	12300	)	,
(	12297	)	,
(	12294	)	,
(	12291	)	,
(	12288	)	,
(	12285	)	,
(	12282	)	,
(	12279	)	,
(	12276	)	,
(	12273	)	,
(	12270	)	,
(	12267	)	,
(	12264	)	,
(	12261	)	,
(	12258	)	,
(	12255	)	,
(	12252	)	,
(	12249	)	,
(	12246	)	,
(	12243	)	,
(	12240	)	,
(	12237	)	,
(	12234	)	,
(	12231	)	,
(	12228	)	,
(	12225	)	,
(	12222	)	,
(	12219	)	,
(	12216	)	,
(	12213	)	,
(	12210	)	,
(	12207	)	,
(	12204	)	,
(	12201	)	,
(	12198	)	,
(	12195	)	,
(	12192	)	,
(	12189	)	,
(	12186	)	,
(	12183	)	,
(	12180	)	,
(	12177	)	,
(	12174	)	,
(	12171	)	,
(	12168	)	,
(	12165	)	,
(	12162	)	,
(	12159	)	,
(	12156	)	,
(	12153	)	,
(	12150	)	,
(	12147	)	,
(	12144	)	,
(	12141	)	,
(	12138	)	,
(	12135	)	,
(	12132	)	,
(	12129	)	,
(	12126	)	,
(	12123	)	,
(	12120	)	,
(	12117	)	,
(	12114	)	,
(	12111	)	,
(	12108	)	,
(	12105	)	,
(	12102	)	,
(	12099	)	,
(	12096	)	,
(	12093	)	,
(	12090	)	,
(	12087	)	,
(	12084	)	,
(	12081	)	,
(	12078	)	,
(	12075	)	,
(	12072	)	,
(	12069	)	,
(	12066	)	,
(	12063	)	,
(	12060	)	,
(	12057	)	,
(	12054	)	,
(	12051	)	,
(	12048	)	,
(	12045	)	,
(	12042	)	,
(	12039	)	,
(	12036	)	,
(	12033	)	,
(	12030	)	,
(	12027	)	,
(	12024	)	,
(	12021	)	,
(	12018	)	,
(	12015	)	,
(	12012	)	,
(	12009	)	,
(	12006	)	,
(	12003	)	,
(	12000	)	,
(	11997	)	,
(	11994	)	,
(	11991	)	,
(	11988	)	,
(	11985	)	,
(	11982	)	,
(	11979	)	,
(	11976	)	,
(	11973	)	,
(	11970	)	,
(	11967	)	,
(	11964	)	,
(	11961	)	,
(	11958	)	,
(	11955	)	,
(	11952	)	,
(	11949	)	,
(	11946	)	,
(	11943	)	,
(	11940	)	,
(	11937	)	,
(	11934	)	,
(	11931	)	,
(	11928	)	,
(	11925	)	,
(	11922	)	,
(	11919	)	,
(	11916	)	,
(	11913	)	,
(	11910	)	,
(	11907	)	,
(	11904	)	,
(	11901	)	,
(	11898	)	,
(	11895	)	,
(	11892	)	,
(	11889	)	,
(	11886	)	,
(	11883	)	,
(	11880	)	,
(	11877	)	,
(	11874	)	,
(	11871	)	,
(	11868	)	,
(	11865	)	,
(	11862	)	,
(	11859	)	,
(	11856	)	,
(	11853	)	,
(	11850	)	,
(	11847	)	,
(	11844	)	,
(	11841	)	,
(	11838	)	,
(	11835	)	,
(	11832	)	,
(	11829	)	,
(	11826	)	,
(	11823	)	,
(	11820	)	,
(	11817	)	,
(	11814	)	,
(	11811	)	,
(	11808	)	,
(	11805	)	,
(	11802	)	,
(	11799	)	,
(	11796	)	,
(	11793	)	,
(	11790	)	,
(	11787	)	,
(	11784	)	,
(	11781	)	,
(	11778	)	,
(	11775	)	,
(	11772	)	,
(	11769	)	,
(	11766	)	,
(	11763	)	,
(	11760	)	,
(	11757	)	,
(	11754	)	,
(	11751	)	,
(	11748	)	,
(	11745	)	,
(	11742	)	,
(	11739	)	,
(	11736	)	,
(	11733	)	,
(	11730	)	,
(	11727	)	,
(	11724	)	,
(	11721	)	,
(	11718	)	,
(	11715	)	,
(	11712	)	,
(	11709	)	,
(	11706	)	,
(	11703	)	,
(	11700	)	,
(	11697	)	,
(	11694	)	,
(	11691	)	,
(	11688	)	,
(	11685	)	,
(	11682	)	,
(	11679	)	,
(	11676	)	,
(	11673	)	,
(	11670	)	,
(	11667	)	,
(	11664	)	,
(	11661	)	,
(	11658	)	,
(	11655	)	,
(	11652	)	,
(	11649	)	,
(	11646	)	,
(	11643	)	,
(	11640	)	,
(	11637	)	,
(	11634	)	,
(	11631	)	,
(	11628	)	,
(	11625	)	,
(	11622	)	,
(	11619	)	,
(	11616	)	,
(	11613	)	,
(	11610	)	,
(	11607	)	,
(	11604	)	,
(	11601	)	,
(	11598	)	,
(	11595	)	,
(	11592	)	,
(	11589	)	,
(	11586	)	,
(	11583	)	,
(	11580	)	,
(	11577	)	,
(	11574	)	,
(	11571	)	,
(	11568	)	,
(	11565	)	,
(	11562	)	,
(	11559	)	,
(	11556	)	,
(	11553	)	,
(	11550	)	,
(	11547	)	,
(	11544	)	,
(	11541	)	,
(	11538	)	,
(	11535	)	,
(	11532	)	,
(	11529	)	,
(	11526	)	,
(	11523	)	,
(	11520	)	,
(	11517	)	,
(	11514	)	,
(	11511	)	,
(	11508	)	,
(	11505	)	,
(	11502	)	,
(	11499	)	,
(	11496	)	,
(	11493	)	,
(	11490	)	,
(	11487	)	,
(	11484	)	,
(	11481	)	,
(	11478	)	,
(	11475	)	,
(	11472	)	,
(	11469	)	,
(	11466	)	,
(	11463	)	,
(	11460	)	,
(	11457	)	,
(	11454	)	,
(	11451	)	,
(	11448	)	,
(	11445	)	,
(	11442	)	,
(	11439	)	,
(	11436	)	,
(	11433	)	,
(	11430	)	,
(	11427	)	,
(	11424	)	,
(	11421	)	,
(	11418	)	,
(	11415	)	,
(	11412	)	,
(	11409	)	,
(	11406	)	,
(	11403	)	,
(	11400	)	,
(	11397	)	,
(	11394	)	,
(	11391	)	,
(	11388	)	,
(	11385	)	,
(	11382	)	,
(	11379	)	,
(	11376	)	,
(	11373	)	,
(	11370	)	,
(	11367	)	,
(	11364	)	,
(	11361	)	,
(	11358	)	,
(	11355	)	,
(	11352	)	,
(	11349	)	,
(	11346	)	,
(	11343	)	,
(	11340	)	,
(	11337	)	,
(	11334	)	,
(	11331	)	,
(	11328	)	,
(	11325	)	,
(	11322	)	,
(	11319	)	,
(	11316	)	,
(	11313	)	,
(	11310	)	,
(	11307	)	,
(	11304	)	,
(	11301	)	,
(	11298	)	,
(	11295	)	,
(	11292	)	,
(	11289	)	,
(	11286	)	,
(	11283	)	,
(	11280	)	,
(	11277	)	,
(	11274	)	,
(	11271	)	,
(	11268	)	,
(	11265	)	,
(	11262	)	,
(	11259	)	,
(	11256	)	,
(	11253	)	,
(	11250	)	,
(	11247	)	,
(	11244	)	,
(	11241	)	,
(	11238	)	,
(	11235	)	,
(	11232	)	,
(	11229	)	,
(	11226	)	,
(	11223	)	,
(	11220	)	,
(	11217	)	,
(	11214	)	,
(	11211	)	,
(	11208	)	,
(	11205	)	,
(	11202	)	,
(	11199	)	,
(	11196	)	,
(	11193	)	,
(	11190	)	,
(	11187	)	,
(	11184	)	,
(	11181	)	,
(	11178	)	,
(	11175	)	,
(	11172	)	,
(	11169	)	,
(	11166	)	,
(	11163	)	,
(	11160	)	,
(	11157	)	,
(	11154	)	,
(	11151	)	,
(	11148	)	,
(	11145	)	,
(	11142	)	,
(	11139	)	,
(	11136	)	,
(	11133	)	,
(	11130	)	,
(	11127	)	,
(	11124	)	,
(	11121	)	,
(	11118	)	,
(	11115	)	,
(	11112	)	,
(	11109	)	,
(	11106	)	,
(	11103	)	,
(	11100	)	,
(	11097	)	,
(	11094	)	,
(	11091	)	,
(	11088	)	,
(	11085	)	,
(	11082	)	,
(	11079	)	,
(	11076	)	,
(	11073	)	,
(	11070	)	,
(	11067	)	,
(	11064	)	,
(	11061	)	,
(	11058	)	,
(	11055	)	,
(	11052	)	,
(	11049	)	,
(	11046	)	,
(	11043	)	,
(	11040	)	,
(	11037	)	,
(	11034	)	,
(	11031	)	,
(	11028	)	,
(	11025	)	,
(	11022	)	,
(	11019	)	,
(	11016	)	,
(	11013	)	,
(	11010	)	,
(	11007	)	,
(	11004	)	,
(	11001	)	,
(	10998	)	,
(	10995	)	,
(	10992	)	,
(	10989	)	,
(	10986	)	,
(	10983	)	,
(	10980	)	,
(	10977	)	,
(	10974	)	,
(	10971	)	,
(	10968	)	,
(	10965	)	,
(	10962	)	,
(	10959	)	,
(	10956	)	,
(	10953	)	,
(	10950	)	,
(	10947	)	,
(	10944	)	,
(	10941	)	,
(	10938	)	,
(	10935	)	,
(	10932	)	,
(	10929	)	,
(	10926	)	,
(	10923	)	,
(	10920	)	,
(	10917	)	,
(	10914	)	,
(	10911	)	,
(	10908	)	,
(	10905	)	,
(	10902	)	,
(	10899	)	,
(	10896	)	,
(	10893	)	,
(	10890	)	,
(	10887	)	,
(	10884	)	,
(	10881	)	,
(	10878	)	,
(	10875	)	,
(	10872	)	,
(	10869	)	,
(	10866	)	,
(	10863	)	,
(	10860	)	,
(	10857	)	,
(	10854	)	,
(	10851	)	,
(	10848	)	,
(	10845	)	,
(	10842	)	,
(	10839	)	,
(	10836	)	,
(	10833	)	,
(	10830	)	,
(	10827	)	,
(	10824	)	,
(	10821	)	,
(	10818	)	,
(	10815	)	,
(	10812	)	,
(	10809	)	,
(	10806	)	,
(	10803	)	,
(	10800	)	,
(	10797	)	,
(	10794	)	,
(	10791	)	,
(	10788	)	,
(	10785	)	,
(	10782	)	,
(	10779	)	,
(	10776	)	,
(	10773	)	,
(	10770	)	,
(	10767	)	,
(	10764	)	,
(	10761	)	,
(	10758	)	,
(	10755	)	,
(	10752	)	,
(	10749	)	,
(	10746	)	,
(	10743	)	,
(	10740	)	,
(	10737	)	,
(	10734	)	,
(	10731	)	,
(	10728	)	,
(	10725	)	,
(	10722	)	,
(	10719	)	,
(	10716	)	,
(	10713	)	,
(	10710	)	,
(	10707	)	,
(	10704	)	,
(	10701	)	,
(	10698	)	,
(	10695	)	,
(	10692	)	,
(	10689	)	,
(	10686	)	,
(	10683	)	,
(	10680	)	,
(	10677	)	,
(	10674	)	,
(	10671	)	,
(	10668	)	,
(	10665	)	,
(	10662	)	,
(	10659	)	,
(	10656	)	,
(	10653	)	,
(	10650	)	,
(	10647	)	,
(	10644	)	,
(	10641	)	,
(	10638	)	,
(	10635	)	,
(	10632	)	,
(	10629	)	,
(	10626	)	,
(	10623	)	,
(	10620	)	,
(	10617	)	,
(	10614	)	,
(	10611	)	,
(	10608	)	,
(	10605	)	,
(	10602	)	,
(	10599	)	,
(	10596	)	,
(	10593	)	,
(	10590	)	,
(	10587	)	,
(	10584	)	,
(	10581	)	,
(	10578	)	,
(	10575	)	,
(	10572	)	,
(	10569	)	,
(	10566	)	,
(	10563	)	,
(	10560	)	,
(	10557	)	,
(	10554	)	,
(	10551	)	,
(	10548	)	,
(	10545	)	,
(	10542	)	,
(	10539	)	,
(	10536	)	,
(	10533	)	,
(	10530	)	,
(	10527	)	,
(	10524	)	,
(	10521	)	,
(	10518	)	,
(	10515	)	,
(	10512	)	,
(	10509	)	,
(	10506	)	,
(	10503	)	,
(	10500	)	,
(	10497	)	,
(	10494	)	,
(	10491	)	,
(	10488	)	,
(	10485	)	,
(	10482	)	,
(	10479	)	,
(	10476	)	,
(	10473	)	,
(	10470	)	,
(	10467	)	,
(	10464	)	,
(	10461	)	,
(	10458	)	,
(	10455	)	,
(	10452	)	,
(	10449	)	,
(	10446	)	,
(	10443	)	,
(	10440	)	,
(	10437	)	,
(	10434	)	,
(	10431	)	,
(	10428	)	,
(	10425	)	,
(	10422	)	,
(	10419	)	,
(	10416	)	,
(	10413	)	,
(	10410	)	,
(	10407	)	,
(	10404	)	,
(	10401	)	,
(	10398	)	,
(	10395	)	,
(	10392	)	,
(	10389	)	,
(	10386	)	,
(	10383	)	,
(	10380	)	,
(	10377	)	,
(	10374	)	,
(	10371	)	,
(	10368	)	,
(	10365	)	,
(	10362	)	,
(	10359	)	,
(	10356	)	,
(	10353	)	,
(	10350	)	,
(	10347	)	,
(	10344	)	,
(	10341	)	,
(	10338	)	,
(	10335	)	,
(	10332	)	,
(	10329	)	,
(	10326	)	,
(	10323	)	,
(	10320	)	,
(	10317	)	,
(	10314	)	,
(	10311	)	,
(	10308	)	,
(	10305	)	,
(	10302	)	,
(	10299	)	,
(	10296	)	,
(	10293	)	,
(	10290	)	,
(	10287	)	,
(	10284	)	,
(	10281	)	,
(	10278	)	,
(	10275	)	,
(	10272	)	,
(	10269	)	,
(	10266	)	,
(	10263	)	,
(	10260	)	,
(	10257	)	,
(	10254	)	,
(	10251	)	,
(	10248	)	,
(	10245	)	,
(	10242	)	,
(	10239	)	,
(	10236	)	,
(	10233	)	,
(	10230	)	,
(	10227	)	,
(	10224	)	,
(	10221	)	,
(	10218	)	,
(	10215	)	,
(	10212	)	,
(	10209	)	,
(	10206	)	,
(	10203	)	,
(	10200	)	,
(	10197	)	,
(	10194	)	,
(	10191	)	,
(	10188	)	,
(	10185	)	,
(	10182	)	,
(	10179	)	,
(	10176	)	,
(	10173	)	,
(	10170	)	,
(	10167	)	,
(	10164	)	,
(	10161	)	,
(	10158	)	,
(	10155	)	,
(	10152	)	,
(	10149	)	,
(	10146	)	,
(	10143	)	,
(	10140	)	,
(	10137	)	,
(	10134	)	,
(	10131	)	,
(	10128	)	,
(	10125	)	,
(	10122	)	,
(	10119	)	,
(	10116	)	,
(	10113	)	,
(	10110	)	,
(	10107	)	,
(	10104	)	,
(	10101	)	,
(	10098	)	,
(	10095	)	,
(	10092	)	,
(	10089	)	,
(	10086	)	,
(	10083	)	,
(	10080	)	,
(	10077	)	,
(	10074	)	,
(	10071	)	,
(	10068	)	,
(	10065	)	,
(	10062	)	,
(	10059	)	,
(	10056	)	,
(	10053	)	,
(	10050	)	,
(	10047	)	,
(	10044	)	,
(	10041	)	,
(	10038	)	,
(	10035	)	,
(	10032	)	,
(	10029	)	,
(	10026	)	,
(	10023	)	,
(	10020	)	,
(	10017	)	,
(	10014	)	,
(	10011	)	,
(	10008	)	,
(	10005	)	,
(	10002	)	,
(	9999	)	,
(	9996	)	,
(	9993	)	,
(	9990	)	,
(	9987	)	,
(	9984	)	,
(	9981	)	,
(	9978	)	,
(	9975	)	,
(	9972	)	,
(	9969	)	,
(	9966	)	,
(	9963	)	,
(	9960	)	,
(	9957	)	,
(	9954	)	,
(	9951	)	,
(	9948	)	,
(	9945	)	,
(	9942	)	,
(	9939	)	,
(	9936	)	,
(	9933	)	,
(	9930	)	,
(	9927	)	,
(	9924	)	,
(	9921	)	,
(	9918	)	,
(	9915	)	,
(	9912	)	,
(	9909	)	,
(	9906	)	,
(	9903	)	,
(	9900	)	,
(	9897	)	,
(	9894	)	,
(	9891	)	,
(	9888	)	,
(	9885	)	,
(	9882	)	,
(	9879	)	,
(	9876	)	,
(	9873	)	,
(	9870	)	,
(	9867	)	,
(	9864	)	,
(	9861	)	,
(	9858	)	,
(	9855	)	,
(	9852	)	,
(	9849	)	,
(	9846	)	,
(	9843	)	,
(	9840	)	,
(	9837	)	,
(	9834	)	,
(	9831	)	,
(	9828	)	,
(	9825	)	,
(	9822	)	,
(	9819	)	,
(	9816	)	,
(	9813	)	,
(	9810	)	,
(	9807	)	,
(	9804	)	,
(	9801	)	,
(	9798	)	,
(	9795	)	,
(	9792	)	,
(	9789	)	,
(	9786	)	,
(	9783	)	,
(	9780	)	,
(	9777	)	,
(	9774	)	,
(	9771	)	,
(	9768	)	,
(	9765	)	,
(	9762	)	,
(	9759	)	,
(	9756	)	,
(	9753	)	,
(	9750	)	,
(	9747	)	,
(	9744	)	,
(	9741	)	,
(	9738	)	,
(	9735	)	,
(	9732	)	,
(	9729	)	,
(	9726	)	,
(	9723	)	,
(	9720	)	,
(	9717	)	,
(	9714	)	,
(	9711	)	,
(	9708	)	,
(	9705	)	,
(	9702	)	,
(	9699	)	,
(	9696	)	,
(	9693	)	,
(	9690	)	,
(	9687	)	,
(	9684	)	,
(	9681	)	,
(	9678	)	,
(	9675	)	,
(	9672	)	,
(	9669	)	,
(	9666	)	,
(	9663	)	,
(	9660	)	,
(	9657	)	,
(	9654	)	,
(	9651	)	,
(	9648	)	,
(	9645	)	,
(	9642	)	,
(	9639	)	,
(	9636	)	,
(	9633	)	,
(	9630	)	,
(	9627	)	,
(	9624	)	,
(	9621	)	,
(	9618	)	,
(	9615	)	,
(	9612	)	,
(	9609	)	,
(	9606	)	,
(	9603	)	,
(	9600	)	,
(	9597	)	,
(	9594	)	,
(	9591	)	,
(	9588	)	,
(	9585	)	,
(	9582	)	,
(	9579	)	,
(	9576	)	,
(	9573	)	,
(	9570	)	,
(	9567	)	,
(	9564	)	,
(	9561	)	,
(	9558	)	,
(	9555	)	,
(	9552	)	,
(	9549	)	,
(	9546	)	,
(	9543	)	,
(	9540	)	,
(	9537	)	,
(	9534	)	,
(	9531	)	,
(	9528	)	,
(	9525	)	,
(	9522	)	,
(	9519	)	,
(	9516	)	,
(	9513	)	,
(	9510	)	,
(	9507	)	,
(	9504	)	,
(	9501	)	,
(	9498	)	,
(	9495	)	,
(	9492	)	,
(	9489	)	,
(	9486	)	,
(	9483	)	,
(	9480	)	,
(	9477	)	,
(	9474	)	,
(	9471	)	,
(	9468	)	,
(	9465	)	,
(	9462	)	,
(	9459	)	,
(	9456	)	,
(	9453	)	,
(	9450	)	,
(	9447	)	,
(	9444	)	,
(	9441	)	,
(	9438	)	,
(	9435	)	,
(	9432	)	,
(	9429	)	,
(	9426	)	,
(	9423	)	,
(	9420	)	,
(	9417	)	,
(	9414	)	,
(	9411	)	,
(	9408	)	,
(	9405	)	,
(	9402	)	,
(	9399	)	,
(	9396	)	,
(	9393	)	,
(	9390	)	,
(	9387	)	,
(	9384	)	,
(	9381	)	,
(	9378	)	,
(	9375	)	,
(	9372	)	,
(	9369	)	,
(	9366	)	,
(	9363	)	,
(	9360	)	,
(	9357	)	,
(	9354	)	,
(	9351	)	,
(	9348	)	,
(	9345	)	,
(	9342	)	,
(	9339	)	,
(	9336	)	,
(	9333	)	,
(	9330	)	,
(	9327	)	,
(	9324	)	,
(	9321	)	,
(	9318	)	,
(	9315	)	,
(	9312	)	,
(	9309	)	,
(	9306	)	,
(	9303	)	,
(	9300	)	,
(	9297	)	,
(	9294	)	,
(	9291	)	,
(	9288	)	,
(	9285	)	,
(	9282	)	,
(	9279	)	,
(	9276	)	,
(	9273	)	,
(	9270	)	,
(	9267	)	,
(	9264	)	,
(	9261	)	,
(	9258	)	,
(	9255	)	,
(	9252	)	,
(	9249	)	,
(	9246	)	,
(	9243	)	,
(	9240	)	,
(	9237	)	,
(	9234	)	,
(	9231	)	,
(	9228	)	,
(	9225	)	,
(	9222	)	,
(	9219	)	,
(	9216	)	,
(	9213	)	,
(	9210	)	,
(	9207	)	,
(	9204	)	,
(	9201	)	,
(	9198	)	,
(	9195	)	,
(	9192	)	,
(	9189	)	,
(	9186	)	,
(	9183	)	,
(	9180	)	,
(	9177	)	,
(	9174	)	,
(	9171	)	,
(	9168	)	,
(	9165	)	,
(	9162	)	,
(	9159	)	,
(	9156	)	,
(	9153	)	,
(	9150	)	,
(	9147	)	,
(	9144	)	,
(	9141	)	,
(	9138	)	,
(	9135	)	,
(	9132	)	,
(	9129	)	,
(	9126	)	,
(	9123	)	,
(	9120	)	,
(	9117	)	,
(	9114	)	,
(	9111	)	,
(	9108	)	,
(	9105	)	,
(	9102	)	,
(	9099	)	,
(	9096	)	,
(	9093	)	,
(	9090	)	,
(	9087	)	,
(	9084	)	,
(	9081	)	,
(	9078	)	,
(	9075	)	,
(	9072	)	,
(	9069	)	,
(	9066	)	,
(	9063	)	,
(	9060	)	,
(	9057	)	,
(	9054	)	,
(	9051	)	,
(	9048	)	,
(	9045	)	,
(	9042	)	,
(	9039	)	,
(	9036	)	,
(	9033	)	,
(	9030	)	,
(	9027	)	,
(	9024	)	,
(	9021	)	,
(	9018	)	,
(	9015	)	,
(	9012	)	,
(	9009	)	,
(	9006	)	,
(	9003	)	,
(	9000	)	,
(	8997	)	,
(	8994	)	,
(	8991	)	,
(	8988	)	,
(	8985	)	,
(	8982	)	,
(	8979	)	,
(	8976	)	,
(	8973	)	,
(	8970	)	,
(	8967	)	,
(	8964	)	,
(	8961	)	,
(	8958	)	,
(	8955	)	,
(	8952	)	,
(	8949	)	,
(	8946	)	,
(	8943	)	,
(	8940	)	,
(	8937	)	,
(	8934	)	,
(	8931	)	,
(	8928	)	,
(	8925	)	,
(	8922	)	,
(	8919	)	,
(	8916	)	,
(	8913	)	,
(	8910	)	,
(	8907	)	,
(	8904	)	,
(	8901	)	,
(	8898	)	,
(	8895	)	,
(	8892	)	,
(	8889	)	,
(	8886	)	,
(	8883	)	,
(	8880	)	,
(	8877	)	,
(	8874	)	,
(	8871	)	,
(	8868	)	,
(	8865	)	,
(	8862	)	,
(	8859	)	,
(	8856	)	,
(	8853	)	,
(	8850	)	,
(	8847	)	,
(	8844	)	,
(	8841	)	,
(	8838	)	,
(	8835	)	,
(	8832	)	,
(	8829	)	,
(	8826	)	,
(	8823	)	,
(	8820	)	,
(	8817	)	,
(	8814	)	,
(	8811	)	,
(	8808	)	,
(	8805	)	,
(	8802	)	,
(	8799	)	,
(	8796	)	,
(	8793	)	,
(	8790	)	,
(	8787	)	,
(	8784	)	,
(	8781	)	,
(	8778	)	,
(	8775	)	,
(	8772	)	,
(	8769	)	,
(	8766	)	,
(	8763	)	,
(	8760	)	,
(	8757	)	,
(	8754	)	,
(	8751	)	,
(	8748	)	,
(	8745	)	,
(	8742	)	,
(	8739	)	,
(	8736	)	,
(	8733	)	,
(	8730	)	,
(	8727	)	,
(	8724	)	,
(	8721	)	,
(	8718	)	,
(	8715	)	,
(	8712	)	,
(	8709	)	,
(	8706	)	,
(	8703	)	,
(	8700	)	,
(	8697	)	,
(	8694	)	,
(	8691	)	,
(	8688	)	,
(	8685	)	,
(	8682	)	,
(	8679	)	,
(	8676	)	,
(	8673	)	,
(	8670	)	,
(	8667	)	,
(	8664	)	,
(	8661	)	,
(	8658	)	,
(	8655	)	,
(	8652	)	,
(	8649	)	,
(	8646	)	,
(	8643	)	,
(	8640	)	,
(	8637	)	,
(	8634	)	,
(	8631	)	,
(	8628	)	,
(	8625	)	,
(	8622	)	,
(	8619	)	,
(	8616	)	,
(	8613	)	,
(	8610	)	,
(	8607	)	,
(	8604	)	,
(	8601	)	,
(	8598	)	,
(	8595	)	,
(	8592	)	,
(	8589	)	,
(	8586	)	,
(	8583	)	,
(	8580	)	,
(	8577	)	,
(	8574	)	,
(	8571	)	,
(	8568	)	,
(	8565	)	,
(	8562	)	,
(	8559	)	,
(	8556	)	,
(	8553	)	,
(	8550	)	,
(	8547	)	,
(	8544	)	,
(	8541	)	,
(	8538	)	,
(	8535	)	,
(	8532	)	,
(	8529	)	,
(	8526	)	,
(	8523	)	,
(	8520	)	,
(	8517	)	,
(	8514	)	,
(	8511	)	,
(	8508	)	,
(	8505	)	,
(	8502	)	,
(	8499	)	,
(	8496	)	,
(	8493	)	,
(	8490	)	,
(	8487	)	,
(	8484	)	,
(	8481	)	,
(	8478	)	,
(	8475	)	,
(	8472	)	,
(	8469	)	,
(	8466	)	,
(	8463	)	,
(	8460	)	,
(	8457	)	,
(	8454	)	,
(	8451	)	,
(	8448	)	,
(	8445	)	,
(	8442	)	,
(	8439	)	,
(	8436	)	,
(	8433	)	,
(	8430	)	,
(	8427	)	,
(	8424	)	,
(	8421	)	,
(	8418	)	,
(	8415	)	,
(	8412	)	,
(	8409	)	,
(	8406	)	,
(	8403	)	,
(	8400	)	,
(	8397	)	,
(	8394	)	,
(	8391	)	,
(	8388	)	,
(	8385	)	,
(	8382	)	,
(	8379	)	,
(	8376	)	,
(	8373	)	,
(	8370	)	,
(	8367	)	,
(	8364	)	,
(	8361	)	,
(	8358	)	,
(	8355	)	,
(	8352	)	,
(	8349	)	,
(	8346	)	,
(	8343	)	,
(	8340	)	,
(	8337	)	,
(	8334	)	,
(	8331	)	,
(	8328	)	,
(	8325	)	,
(	8322	)	,
(	8319	)	,
(	8316	)	,
(	8313	)	,
(	8310	)	,
(	8307	)	,
(	8304	)	,
(	8301	)	,
(	8298	)	,
(	8295	)	,
(	8292	)	,
(	8289	)	,
(	8286	)	,
(	8283	)	,
(	8280	)	,
(	8277	)	,
(	8274	)	,
(	8271	)	,
(	8268	)	,
(	8265	)	,
(	8262	)	,
(	8259	)	,
(	8256	)	,
(	8253	)	,
(	8250	)	,
(	8247	)	,
(	8244	)	,
(	8241	)	,
(	8238	)	,
(	8235	)	,
(	8232	)	,
(	8229	)	,
(	8226	)	,
(	8223	)	,
(	8220	)	,
(	8217	)	,
(	8214	)	,
(	8211	)	,
(	8208	)	,
(	8205	)	,
(	8202	)	,
(	8199	)	,
(	8196	)	,
(	8193	)	,
(	8190	)	,
(	8187	)	,
(	8184	)	,
(	8181	)	,
(	8178	)	,
(	8175	)	,
(	8172	)	,
(	8169	)	,
(	8166	)	,
(	8163	)	,
(	8160	)	,
(	8157	)	,
(	8154	)	,
(	8151	)	,
(	8148	)	,
(	8145	)	,
(	8142	)	,
(	8139	)	,
(	8136	)	,
(	8133	)	,
(	8130	)	,
(	8127	)	,
(	8124	)	,
(	8121	)	,
(	8118	)	,
(	8115	)	,
(	8112	)	,
(	8109	)	,
(	8106	)	,
(	8103	)	,
(	8100	)	,
(	8097	)	,
(	8094	)	,
(	8091	)	,
(	8088	)	,
(	8085	)	,
(	8082	)	,
(	8079	)	,
(	8076	)	,
(	8073	)	,
(	8070	)	,
(	8067	)	,
(	8064	)	,
(	8061	)	,
(	8058	)	,
(	8055	)	,
(	8052	)	,
(	8049	)	,
(	8046	)	,
(	8043	)	,
(	8040	)	,
(	8037	)	,
(	8034	)	,
(	8031	)	,
(	8028	)	,
(	8025	)	,
(	8022	)	,
(	8019	)	,
(	8016	)	,
(	8013	)	,
(	8010	)	,
(	8007	)	,
(	8004	)	,
(	8001	)	,
(	7998	)	,
(	7995	)	,
(	7992	)	,
(	7989	)	,
(	7986	)	,
(	7983	)	,
(	7980	)	,
(	7977	)	,
(	7974	)	,
(	7971	)	,
(	7968	)	,
(	7965	)	,
(	7962	)	,
(	7959	)	,
(	7956	)	,
(	7953	)	,
(	7950	)	,
(	7947	)	,
(	7944	)	,
(	7941	)	,
(	7938	)	,
(	7935	)	,
(	7932	)	,
(	7929	)	,
(	7926	)	,
(	7923	)	,
(	7920	)	,
(	7917	)	,
(	7914	)	,
(	7911	)	,
(	7908	)	,
(	7905	)	,
(	7902	)	,
(	7899	)	,
(	7896	)	,
(	7893	)	,
(	7890	)	,
(	7887	)	,
(	7884	)	,
(	7881	)	,
(	7878	)	,
(	7875	)	,
(	7872	)	,
(	7869	)	,
(	7866	)	,
(	7863	)	,
(	7860	)	,
(	7857	)	,
(	7854	)	,
(	7851	)	,
(	7848	)	,
(	7845	)	,
(	7842	)	,
(	7839	)	,
(	7836	)	,
(	7833	)	,
(	7830	)	,
(	7827	)	,
(	7824	)	,
(	7821	)	,
(	7818	)	,
(	7815	)	,
(	7812	)	,
(	7809	)	,
(	7806	)	,
(	7803	)	,
(	7800	)	,
(	7797	)	,
(	7794	)	,
(	7791	)	,
(	7788	)	,
(	7785	)	,
(	7782	)	,
(	7779	)	,
(	7776	)	,
(	7773	)	,
(	7770	)	,
(	7767	)	,
(	7764	)	,
(	7761	)	,
(	7758	)	,
(	7755	)	,
(	7752	)	,
(	7749	)	,
(	7746	)	,
(	7743	)	,
(	7740	)	,
(	7737	)	,
(	7734	)	,
(	7731	)	,
(	7728	)	,
(	7725	)	,
(	7722	)	,
(	7719	)	,
(	7716	)	,
(	7713	)	,
(	7710	)	,
(	7707	)	,
(	7704	)	,
(	7701	)	,
(	7698	)	,
(	7695	)	,
(	7692	)	,
(	7689	)	,
(	7686	)	,
(	7683	)	,
(	7680	)	,
(	7677	)	,
(	7674	)	,
(	7671	)	,
(	7668	)	,
(	7665	)	,
(	7662	)	,
(	7659	)	,
(	7656	)	,
(	7653	)	,
(	7650	)	,
(	7647	)	,
(	7644	)	,
(	7641	)	,
(	7638	)	,
(	7635	)	,
(	7632	)	,
(	7629	)	,
(	7626	)	,
(	7623	)	,
(	7620	)	,
(	7617	)	,
(	7614	)	,
(	7611	)	,
(	7608	)	,
(	7605	)	,
(	7602	)	,
(	7599	)	,
(	7596	)	,
(	7593	)	,
(	7590	)	,
(	7587	)	,
(	7584	)	,
(	7581	)	,
(	7578	)	,
(	7575	)	,
(	7572	)	,
(	7569	)	,
(	7566	)	,
(	7563	)	,
(	7560	)	,
(	7557	)	,
(	7554	)	,
(	7551	)	,
(	7548	)	,
(	7545	)	,
(	7542	)	,
(	7539	)	,
(	7536	)	,
(	7533	)	,
(	7530	)	,
(	7527	)	,
(	7524	)	,
(	7521	)	,
(	7518	)	,
(	7515	)	,
(	7512	)	,
(	7509	)	,
(	7506	)	,
(	7503	)	,
(	7500	)	,
(	7497	)	,
(	7494	)	,
(	7491	)	,
(	7488	)	,
(	7485	)	,
(	7482	)	,
(	7479	)	,
(	7476	)	,
(	7473	)	,
(	7470	)	,
(	7467	)	,
(	7464	)	,
(	7461	)	,
(	7458	)	,
(	7455	)	,
(	7452	)	,
(	7449	)	,
(	7446	)	,
(	7443	)	,
(	7440	)	,
(	7437	)	,
(	7434	)	,
(	7431	)	,
(	7428	)	,
(	7425	)	,
(	7422	)	,
(	7419	)	,
(	7416	)	,
(	7413	)	,
(	7410	)	,
(	7407	)	,
(	7404	)	,
(	7401	)	,
(	7398	)	,
(	7395	)	,
(	7392	)	,
(	7389	)	,
(	7386	)	,
(	7383	)	,
(	7380	)	,
(	7377	)	,
(	7374	)	,
(	7371	)	,
(	7368	)	,
(	7365	)	,
(	7362	)	,
(	7359	)	,
(	7356	)	,
(	7353	)	,
(	7350	)	,
(	7347	)	,
(	7344	)	,
(	7341	)	,
(	7338	)	,
(	7335	)	,
(	7332	)	,
(	7329	)	,
(	7326	)	,
(	7323	)	,
(	7320	)	,
(	7317	)	,
(	7314	)	,
(	7311	)	,
(	7308	)	,
(	7305	)	,
(	7302	)	,
(	7299	)	,
(	7296	)	,
(	7293	)	,
(	7290	)	,
(	7287	)	,
(	7284	)	,
(	7281	)	,
(	7278	)	,
(	7275	)	,
(	7272	)	,
(	7269	)	,
(	7266	)	,
(	7263	)	,
(	7260	)	,
(	7257	)	,
(	7254	)	,
(	7251	)	,
(	7248	)	,
(	7245	)	,
(	7242	)	,
(	7239	)	,
(	7236	)	,
(	7233	)	,
(	7230	)	,
(	7227	)	,
(	7224	)	,
(	7221	)	,
(	7218	)	,
(	7215	)	,
(	7212	)	,
(	7209	)	,
(	7206	)	,
(	7203	)	,
(	7200	)	,
(	7197	)	,
(	7194	)	,
(	7191	)	,
(	7188	)	,
(	7185	)	,
(	7182	)	,
(	7179	)	,
(	7176	)	,
(	7173	)	,
(	7170	)	,
(	7167	)	,
(	7164	)	,
(	7161	)	,
(	7158	)	,
(	7155	)	,
(	7152	)	,
(	7149	)	,
(	7146	)	,
(	7143	)	,
(	7140	)	,
(	7137	)	,
(	7134	)	,
(	7131	)	,
(	7128	)	,
(	7125	)	,
(	7122	)	,
(	7119	)	,
(	7116	)	,
(	7113	)	,
(	7110	)	,
(	7107	)	,
(	7104	)	,
(	7101	)	,
(	7098	)	,
(	7095	)	,
(	7092	)	,
(	7089	)	,
(	7086	)	,
(	7083	)	,
(	7080	)	,
(	7077	)	,
(	7074	)	,
(	7071	)	,
(	7068	)	,
(	7065	)	,
(	7062	)	,
(	7059	)	,
(	7056	)	,
(	7053	)	,
(	7050	)	,
(	7047	)	,
(	7044	)	,
(	7041	)	,
(	7038	)	,
(	7035	)	,
(	7032	)	,
(	7029	)	,
(	7026	)	,
(	7023	)	,
(	7020	)	,
(	7017	)	,
(	7014	)	,
(	7011	)	,
(	7008	)	,
(	7005	)	,
(	7002	)	,
(	6999	)	,
(	6996	)	,
(	6993	)	,
(	6990	)	,
(	6987	)	,
(	6984	)	,
(	6981	)	,
(	6978	)	,
(	6975	)	,
(	6972	)	,
(	6969	)	,
(	6966	)	,
(	6963	)	,
(	6960	)	,
(	6957	)	,
(	6954	)	,
(	6951	)	,
(	6948	)	,
(	6945	)	,
(	6942	)	,
(	6939	)	,
(	6936	)	,
(	6933	)	,
(	6930	)	,
(	6927	)	,
(	6924	)	,
(	6921	)	,
(	6918	)	,
(	6915	)	,
(	6912	)	,
(	6909	)	,
(	6906	)	,
(	6903	)	,
(	6900	)	,
(	6897	)	,
(	6894	)	,
(	6891	)	,
(	6888	)	,
(	6885	)	,
(	6882	)	,
(	6879	)	,
(	6876	)	,
(	6873	)	,
(	6870	)	,
(	6867	)	,
(	6864	)	,
(	6861	)	,
(	6858	)	,
(	6855	)	,
(	6852	)	,
(	6849	)	,
(	6846	)	,
(	6843	)	,
(	6840	)	,
(	6837	)	,
(	6834	)	,
(	6831	)	,
(	6828	)	,
(	6825	)	,
(	6822	)	,
(	6819	)	,
(	6816	)	,
(	6813	)	,
(	6810	)	,
(	6807	)	,
(	6804	)	,
(	6801	)	,
(	6798	)	,
(	6795	)	,
(	6792	)	,
(	6789	)	,
(	6786	)	,
(	6783	)	,
(	6780	)	,
(	6777	)	,
(	6774	)	,
(	6771	)	,
(	6768	)	,
(	6765	)	,
(	6762	)	,
(	6759	)	,
(	6756	)	,
(	6753	)	,
(	6750	)	,
(	6747	)	,
(	6744	)	,
(	6741	)	,
(	6738	)	,
(	6735	)	,
(	6732	)	,
(	6729	)	,
(	6726	)	,
(	6723	)	,
(	6720	)	,
(	6717	)	,
(	6714	)	,
(	6711	)	,
(	6708	)	,
(	6705	)	,
(	6702	)	,
(	6699	)	,
(	6696	)	,
(	6693	)	,
(	6690	)	,
(	6687	)	,
(	6684	)	,
(	6681	)	,
(	6678	)	,
(	6675	)	,
(	6672	)	,
(	6669	)	,
(	6666	)	,
(	6663	)	,
(	6660	)	,
(	6657	)	,
(	6654	)	,
(	6651	)	,
(	6648	)	,
(	6645	)	,
(	6642	)	,
(	6639	)	,
(	6636	)	,
(	6633	)	,
(	6630	)	,
(	6627	)	,
(	6624	)	,
(	6621	)	,
(	6618	)	,
(	6615	)	,
(	6612	)	,
(	6609	)	,
(	6606	)	,
(	6603	)	,
(	6600	)	,
(	6597	)	,
(	6594	)	,
(	6591	)	,
(	6588	)	,
(	6585	)	,
(	6582	)	,
(	6579	)	,
(	6576	)	,
(	6573	)	,
(	6570	)	,
(	6567	)	,
(	6564	)	,
(	6561	)	,
(	6558	)	,
(	6555	)	,
(	6552	)	,
(	6549	)	,
(	6546	)	,
(	6543	)	,
(	6540	)	,
(	6537	)	,
(	6534	)	,
(	6531	)	,
(	6528	)	,
(	6525	)	,
(	6522	)	,
(	6519	)	,
(	6516	)	,
(	6513	)	,
(	6510	)	,
(	6507	)	,
(	6504	)	,
(	6501	)	,
(	6498	)	,
(	6495	)	,
(	6492	)	,
(	6489	)	,
(	6486	)	,
(	6483	)	,
(	6480	)	,
(	6477	)	,
(	6474	)	,
(	6471	)	,
(	6468	)	,
(	6465	)	,
(	6462	)	,
(	6459	)	,
(	6456	)	,
(	6453	)	,
(	6450	)	,
(	6447	)	,
(	6444	)	,
(	6441	)	,
(	6438	)	,
(	6435	)	,
(	6432	)	,
(	6429	)	,
(	6426	)	,
(	6423	)	,
(	6420	)	,
(	6417	)	,
(	6414	)	,
(	6411	)	,
(	6408	)	,
(	6405	)	,
(	6402	)	,
(	6399	)	,
(	6396	)	,
(	6393	)	,
(	6390	)	,
(	6387	)	,
(	6384	)	,
(	6381	)	,
(	6378	)	,
(	6375	)	,
(	6372	)	,
(	6369	)	,
(	6366	)	,
(	6363	)	,
(	6360	)	,
(	6357	)	,
(	6354	)	,
(	6351	)	,
(	6348	)	,
(	6345	)	,
(	6342	)	,
(	6339	)	,
(	6336	)	,
(	6333	)	,
(	6330	)	,
(	6327	)	,
(	6324	)	,
(	6321	)	,
(	6318	)	,
(	6315	)	,
(	6312	)	,
(	6309	)	,
(	6306	)	,
(	6303	)	,
(	6300	)	,
(	6297	)	,
(	6294	)	,
(	6291	)	,
(	6288	)	,
(	6285	)	,
(	6282	)	,
(	6279	)	,
(	6276	)	,
(	6273	)	,
(	6270	)	,
(	6267	)	,
(	6264	)	,
(	6261	)	,
(	6258	)	,
(	6255	)	,
(	6252	)	,
(	6249	)	,
(	6246	)	,
(	6243	)	,
(	6240	)	,
(	6237	)	,
(	6234	)	,
(	6231	)	,
(	6228	)	,
(	6225	)	,
(	6222	)	,
(	6219	)	,
(	6216	)	,
(	6213	)	,
(	6210	)	,
(	6207	)	,
(	6204	)	,
(	6201	)	,
(	6198	)	,
(	6195	)	,
(	6192	)	,
(	6189	)	,
(	6186	)	,
(	6183	)	,
(	6180	)	,
(	6177	)	,
(	6174	)	,
(	6171	)	,
(	6168	)	,
(	6165	)	,
(	6162	)	,
(	6159	)	,
(	6156	)	,
(	6153	)	,
(	6150	)	,
(	6147	)	,
(	6144	)	,
(	6141	)	,
(	6138	)	,
(	6135	)	,
(	6132	)	,
(	6129	)	,
(	6126	)	,
(	6123	)	,
(	6120	)	,
(	6117	)	,
(	6114	)	,
(	6111	)	,
(	6108	)	,
(	6105	)	,
(	6102	)	,
(	6099	)	,
(	6096	)	,
(	6093	)	,
(	6090	)	,
(	6087	)	,
(	6084	)	,
(	6081	)	,
(	6078	)	,
(	6075	)	,
(	6072	)	,
(	6069	)	,
(	6066	)	,
(	6063	)	,
(	6060	)	,
(	6057	)	,
(	6054	)	,
(	6051	)	,
(	6048	)	,
(	6045	)	,
(	6042	)	,
(	6039	)	,
(	6036	)	,
(	6033	)	,
(	6030	)	,
(	6027	)	,
(	6024	)	,
(	6021	)	,
(	6018	)	,
(	6015	)	,
(	6012	)	,
(	6009	)	,
(	6006	)	,
(	6003	)	,
(	6000	)	,
(	5997	)	,
(	5994	)	,
(	5991	)	,
(	5988	)	,
(	5985	)	,
(	5982	)	,
(	5979	)	,
(	5976	)	,
(	5973	)	,
(	5970	)	,
(	5967	)	,
(	5964	)	,
(	5961	)	,
(	5958	)	,
(	5955	)	,
(	5952	)	,
(	5949	)	,
(	5946	)	,
(	5943	)	,
(	5940	)	,
(	5937	)	,
(	5934	)	,
(	5931	)	,
(	5928	)	,
(	5925	)	,
(	5922	)	,
(	5919	)	,
(	5916	)	,
(	5913	)	,
(	5910	)	,
(	5907	)	,
(	5904	)	,
(	5901	)	,
(	5898	)	,
(	5895	)	,
(	5892	)	,
(	5889	)	,
(	5886	)	,
(	5883	)	,
(	5880	)	,
(	5877	)	,
(	5874	)	,
(	5871	)	,
(	5868	)	,
(	5865	)	,
(	5862	)	,
(	5859	)	,
(	5856	)	,
(	5853	)	,
(	5850	)	,
(	5847	)	,
(	5844	)	,
(	5841	)	,
(	5838	)	,
(	5835	)	,
(	5832	)	,
(	5829	)	,
(	5826	)	,
(	5823	)	,
(	5820	)	,
(	5817	)	,
(	5814	)	,
(	5811	)	,
(	5808	)	,
(	5805	)	,
(	5802	)	,
(	5799	)	,
(	5796	)	,
(	5793	)	,
(	5790	)	,
(	5787	)	,
(	5784	)	,
(	5781	)	,
(	5778	)	,
(	5775	)	,
(	5772	)	,
(	5769	)	,
(	5766	)	,
(	5763	)	,
(	5760	)	,
(	5757	)	,
(	5754	)	,
(	5751	)	,
(	5748	)	,
(	5745	)	,
(	5742	)	,
(	5739	)	,
(	5736	)	,
(	5733	)	,
(	5730	)	,
(	5727	)	,
(	5724	)	,
(	5721	)	,
(	5718	)	,
(	5715	)	,
(	5712	)	,
(	5709	)	,
(	5706	)	,
(	5703	)	,
(	5700	)	,
(	5697	)	,
(	5694	)	,
(	5691	)	,
(	5688	)	,
(	5685	)	,
(	5682	)	,
(	5679	)	,
(	5676	)	,
(	5673	)	,
(	5670	)	,
(	5667	)	,
(	5664	)	,
(	5661	)	,
(	5658	)	,
(	5655	)	,
(	5652	)	,
(	5649	)	,
(	5646	)	,
(	5643	)	,
(	5640	)	,
(	5637	)	,
(	5634	)	,
(	5631	)	,
(	5628	)	,
(	5625	)	,
(	5622	)	,
(	5619	)	,
(	5616	)	,
(	5613	)	,
(	5610	)	,
(	5607	)	,
(	5604	)	,
(	5601	)	,
(	5598	)	,
(	5595	)	,
(	5592	)	,
(	5589	)	,
(	5586	)	,
(	5583	)	,
(	5580	)	,
(	5577	)	,
(	5574	)	,
(	5571	)	,
(	5568	)	,
(	5565	)	,
(	5562	)	,
(	5559	)	,
(	5556	)	,
(	5553	)	,
(	5550	)	,
(	5547	)	,
(	5544	)	,
(	5541	)	,
(	5538	)	,
(	5535	)	,
(	5532	)	,
(	5529	)	,
(	5526	)	,
(	5523	)	,
(	5520	)	,
(	5517	)	,
(	5514	)	,
(	5511	)	,
(	5508	)	,
(	5505	)	,
(	5502	)	,
(	5499	)	,
(	5496	)	,
(	5493	)	,
(	5490	)	,
(	5487	)	,
(	5484	)	,
(	5481	)	,
(	5478	)	,
(	5475	)	,
(	5472	)	,
(	5469	)	,
(	5466	)	,
(	5463	)	,
(	5460	)	,
(	5457	)	,
(	5454	)	,
(	5451	)	,
(	5448	)	,
(	5445	)	,
(	5442	)	,
(	5439	)	,
(	5436	)	,
(	5433	)	,
(	5430	)	,
(	5427	)	,
(	5424	)	,
(	5421	)	,
(	5418	)	,
(	5415	)	,
(	5412	)	,
(	5409	)	,
(	5406	)	,
(	5403	)	,
(	5400	)	,
(	5397	)	,
(	5394	)	,
(	5391	)	,
(	5388	)	,
(	5385	)	,
(	5382	)	,
(	5379	)	,
(	5376	)	,
(	5373	)	,
(	5370	)	,
(	5367	)	,
(	5364	)	,
(	5361	)	,
(	5358	)	,
(	5355	)	,
(	5352	)	,
(	5349	)	,
(	5346	)	,
(	5343	)	,
(	5340	)	,
(	5337	)	,
(	5334	)	,
(	5331	)	,
(	5328	)	,
(	5325	)	,
(	5322	)	,
(	5319	)	,
(	5316	)	,
(	5313	)	,
(	5310	)	,
(	5307	)	,
(	5304	)	,
(	5301	)	,
(	5298	)	,
(	5295	)	,
(	5292	)	,
(	5289	)	,
(	5286	)	,
(	5283	)	,
(	5280	)	,
(	5277	)	,
(	5274	)	,
(	5271	)	,
(	5268	)	,
(	5265	)	,
(	5262	)	,
(	5259	)	,
(	5256	)	,
(	5253	)	,
(	5250	)	,
(	5247	)	,
(	5244	)	,
(	5241	)	,
(	5238	)	,
(	5235	)	,
(	5232	)	,
(	5229	)	,
(	5226	)	,
(	5223	)	,
(	5220	)	,
(	5217	)	,
(	5214	)	,
(	5211	)	,
(	5208	)	,
(	5205	)	,
(	5202	)	,
(	5199	)	,
(	5196	)	,
(	5193	)	,
(	5190	)	,
(	5187	)	,
(	5184	)	,
(	5181	)	,
(	5178	)	,
(	5175	)	,
(	5172	)	,
(	5169	)	,
(	5166	)	,
(	5163	)	,
(	5160	)	,
(	5157	)	,
(	5154	)	,
(	5151	)	,
(	5148	)	,
(	5145	)	,
(	5142	)	,
(	5139	)	,
(	5136	)	,
(	5133	)	,
(	5130	)	,
(	5127	)	,
(	5124	)	,
(	5121	)	,
(	5118	)	,
(	5115	)	,
(	5112	)	,
(	5109	)	,
(	5106	)	,
(	5103	)	,
(	5100	)	,
(	5097	)	,
(	5094	)	,
(	5091	)	,
(	5088	)	,
(	5085	)	,
(	5082	)	,
(	5079	)	,
(	5076	)	,
(	5073	)	,
(	5070	)	,
(	5067	)	,
(	5064	)	,
(	5061	)	,
(	5058	)	,
(	5055	)	,
(	5052	)	,
(	5049	)	,
(	5046	)	,
(	5043	)	,
(	5040	)	,
(	5037	)	,
(	5034	)	,
(	5031	)	,
(	5028	)	,
(	5025	)	,
(	5022	)	,
(	5019	)	,
(	5016	)	,
(	5013	)	,
(	5010	)	,
(	5007	)	,
(	5004	)	,
(	5001	)	,
(	4998	)	,
(	4995	)	,
(	4992	)	,
(	4989	)	,
(	4986	)	,
(	4983	)	,
(	4980	)	,
(	4977	)	,
(	4974	)	,
(	4971	)	,
(	4968	)	,
(	4965	)	,
(	4962	)	,
(	4959	)	,
(	4956	)	,
(	4953	)	,
(	4950	)	,
(	4947	)	,
(	4944	)	,
(	4941	)	,
(	4938	)	,
(	4935	)	,
(	4932	)	,
(	4929	)	,
(	4926	)	,
(	4923	)	,
(	4920	)	,
(	4917	)	,
(	4914	)	,
(	4911	)	,
(	4908	)	,
(	4905	)	,
(	4902	)	,
(	4899	)	,
(	4896	)	,
(	4893	)	,
(	4890	)	,
(	4887	)	,
(	4884	)	,
(	4881	)	,
(	4878	)	,
(	4875	)	,
(	4872	)	,
(	4869	)	,
(	4866	)	,
(	4863	)	,
(	4860	)	,
(	4857	)	,
(	4854	)	,
(	4851	)	,
(	4848	)	,
(	4845	)	,
(	4842	)	,
(	4839	)	,
(	4836	)	,
(	4833	)	,
(	4830	)	,
(	4827	)	,
(	4824	)	,
(	4821	)	,
(	4818	)	,
(	4815	)	,
(	4812	)	,
(	4809	)	,
(	4806	)	,
(	4803	)	,
(	4800	)	,
(	4797	)	,
(	4794	)	,
(	4791	)	,
(	4788	)	,
(	4785	)	,
(	4782	)	,
(	4779	)	,
(	4776	)	,
(	4773	)	,
(	4770	)	,
(	4767	)	,
(	4764	)	,
(	4761	)	,
(	4758	)	,
(	4755	)	,
(	4752	)	,
(	4749	)	,
(	4746	)	,
(	4743	)	,
(	4740	)	,
(	4737	)	,
(	4734	)	,
(	4731	)	,
(	4728	)	,
(	4725	)	,
(	4722	)	,
(	4719	)	,
(	4716	)	,
(	4713	)	,
(	4710	)	,
(	4707	)	,
(	4704	)	,
(	4701	)	,
(	4698	)	,
(	4695	)	,
(	4692	)	,
(	4689	)	,
(	4686	)	,
(	4683	)	,
(	4680	)	,
(	4677	)	,
(	4674	)	,
(	4671	)	,
(	4668	)	,
(	4665	)	,
(	4662	)	,
(	4659	)	,
(	4656	)	,
(	4653	)	,
(	4650	)	,
(	4647	)	,
(	4644	)	,
(	4641	)	,
(	4638	)	,
(	4635	)	,
(	4632	)	,
(	4629	)	,
(	4626	)	,
(	4623	)	,
(	4620	)	,
(	4617	)	,
(	4614	)	,
(	4611	)	,
(	4608	)	,
(	4605	)	,
(	4602	)	,
(	4599	)	,
(	4596	)	,
(	4593	)	,
(	4590	)	,
(	4587	)	,
(	4584	)	,
(	4581	)	,
(	4578	)	,
(	4575	)	,
(	4572	)	,
(	4569	)	,
(	4566	)	,
(	4563	)	,
(	4560	)	,
(	4557	)	,
(	4554	)	,
(	4551	)	,
(	4548	)	,
(	4545	)	,
(	4542	)	,
(	4539	)	,
(	4536	)	,
(	4533	)	,
(	4530	)	,
(	4527	)	,
(	4524	)	,
(	4521	)	,
(	4518	)	,
(	4515	)	,
(	4512	)	,
(	4509	)	,
(	4506	)	,
(	4503	)	,
(	4500	)	,
(	4497	)	,
(	4494	)	,
(	4491	)	,
(	4488	)	,
(	4485	)	,
(	4482	)	,
(	4479	)	,
(	4476	)	,
(	4473	)	,
(	4470	)	,
(	4467	)	,
(	4464	)	,
(	4461	)	,
(	4458	)	,
(	4455	)	,
(	4452	)	,
(	4449	)	,
(	4446	)	,
(	4443	)	,
(	4440	)	,
(	4437	)	,
(	4434	)	,
(	4431	)	,
(	4428	)	,
(	4425	)	,
(	4422	)	,
(	4419	)	,
(	4416	)	,
(	4413	)	,
(	4410	)	,
(	4407	)	,
(	4404	)	,
(	4401	)	,
(	4398	)	,
(	4395	)	,
(	4392	)	,
(	4389	)	,
(	4386	)	,
(	4383	)	,
(	4380	)	,
(	4377	)	,
(	4374	)	,
(	4371	)	
 );
 
 end package buzzer_LUT_pkg;