library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4094	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4093	)	,
(	4092	)	,
(	4086	)	,
(	4080	)	,
(	4074	)	,
(	4068	)	,
(	4062	)	,
(	4056	)	,
(	4051	)	,
(	4045	)	,
(	4039	)	,
(	4033	)	,
(	4027	)	,
(	4021	)	,
(	4015	)	,
(	4009	)	,
(	4004	)	,
(	3998	)	,
(	3992	)	,
(	3986	)	,
(	3980	)	,
(	3974	)	,
(	3969	)	,
(	3963	)	,
(	3957	)	,
(	3951	)	,
(	3946	)	,
(	3940	)	,
(	3934	)	,
(	3928	)	,
(	3923	)	,
(	3917	)	,
(	3911	)	,
(	3905	)	,
(	3900	)	,
(	3894	)	,
(	3888	)	,
(	3883	)	,
(	3877	)	,
(	3871	)	,
(	3866	)	,
(	3860	)	,
(	3854	)	,
(	3849	)	,
(	3843	)	,
(	3837	)	,
(	3832	)	,
(	3826	)	,
(	3820	)	,
(	3815	)	,
(	3809	)	,
(	3804	)	,
(	3798	)	,
(	3792	)	,
(	3787	)	,
(	3781	)	,
(	3776	)	,
(	3770	)	,
(	3765	)	,
(	3759	)	,
(	3754	)	,
(	3748	)	,
(	3743	)	,
(	3737	)	,
(	3732	)	,
(	3726	)	,
(	3721	)	,
(	3715	)	,
(	3710	)	,
(	3704	)	,
(	3699	)	,
(	3693	)	,
(	3688	)	,
(	3683	)	,
(	3677	)	,
(	3672	)	,
(	3666	)	,
(	3661	)	,
(	3655	)	,
(	3650	)	,
(	3645	)	,
(	3639	)	,
(	3634	)	,
(	3629	)	,
(	3623	)	,
(	3618	)	,
(	3613	)	,
(	3607	)	,
(	3602	)	,
(	3597	)	,
(	3591	)	,
(	3586	)	,
(	3581	)	,
(	3575	)	,
(	3570	)	,
(	3565	)	,
(	3560	)	,
(	3554	)	,
(	3549	)	,
(	3544	)	,
(	3539	)	,
(	3533	)	,
(	3528	)	,
(	3523	)	,
(	3518	)	,
(	3512	)	,
(	3507	)	,
(	3502	)	,
(	3497	)	,
(	3492	)	,
(	3487	)	,
(	3481	)	,
(	3476	)	,
(	3471	)	,
(	3466	)	,
(	3461	)	,
(	3456	)	,
(	3451	)	,
(	3445	)	,
(	3440	)	,
(	3435	)	,
(	3430	)	,
(	3425	)	,
(	3420	)	,
(	3415	)	,
(	3410	)	,
(	3405	)	,
(	3400	)	,
(	3395	)	,
(	3390	)	,
(	3385	)	,
(	3380	)	,
(	3375	)	,
(	3370	)	,
(	3365	)	,
(	3360	)	,
(	3355	)	,
(	3350	)	,
(	3345	)	,
(	3340	)	,
(	3335	)	,
(	3330	)	,
(	3325	)	,
(	3320	)	,
(	3315	)	,
(	3310	)	,
(	3305	)	,
(	3300	)	,
(	3295	)	,
(	3290	)	,
(	3285	)	,
(	3280	)	,
(	3276	)	,
(	3271	)	,
(	3266	)	,
(	3261	)	,
(	3256	)	,
(	3251	)	,
(	3246	)	,
(	3242	)	,
(	3237	)	,
(	3232	)	,
(	3227	)	,
(	3222	)	,
(	3217	)	,
(	3213	)	,
(	3208	)	,
(	3203	)	,
(	3198	)	,
(	3193	)	,
(	3189	)	,
(	3184	)	,
(	3179	)	,
(	3174	)	,
(	3170	)	,
(	3165	)	,
(	3160	)	,
(	3156	)	,
(	3151	)	,
(	3146	)	,
(	3141	)	,
(	3137	)	,
(	3132	)	,
(	3127	)	,
(	3123	)	,
(	3118	)	,
(	3113	)	,
(	3109	)	,
(	3104	)	,
(	3099	)	,
(	3095	)	,
(	3090	)	,
(	3085	)	,
(	3081	)	,
(	3076	)	,
(	3072	)	,
(	3067	)	,
(	3062	)	,
(	3058	)	,
(	3053	)	,
(	3049	)	,
(	3044	)	,
(	3040	)	,
(	3035	)	,
(	3030	)	,
(	3026	)	,
(	3021	)	,
(	3017	)	,
(	3012	)	,
(	3008	)	,
(	3003	)	,
(	2999	)	,
(	2994	)	,
(	2990	)	,
(	2985	)	,
(	2981	)	,
(	2976	)	,
(	2972	)	,
(	2967	)	,
(	2963	)	,
(	2959	)	,
(	2954	)	,
(	2950	)	,
(	2945	)	,
(	2941	)	,
(	2936	)	,
(	2932	)	,
(	2928	)	,
(	2923	)	,
(	2919	)	,
(	2914	)	,
(	2910	)	,
(	2906	)	,
(	2901	)	,
(	2897	)	,
(	2893	)	,
(	2888	)	,
(	2884	)	,
(	2880	)	,
(	2875	)	,
(	2871	)	,
(	2867	)	,
(	2862	)	,
(	2858	)	,
(	2854	)	,
(	2849	)	,
(	2845	)	,
(	2841	)	,
(	2837	)	,
(	2832	)	,
(	2828	)	,
(	2824	)	,
(	2820	)	,
(	2815	)	,
(	2811	)	,
(	2807	)	,
(	2803	)	,
(	2798	)	,
(	2794	)	,
(	2790	)	,
(	2786	)	,
(	2782	)	,
(	2777	)	,
(	2773	)	,
(	2769	)	,
(	2765	)	,
(	2761	)	,
(	2757	)	,
(	2752	)	,
(	2748	)	,
(	2744	)	,
(	2740	)	,
(	2736	)	,
(	2732	)	,
(	2728	)	,
(	2723	)	,
(	2719	)	,
(	2715	)	,
(	2711	)	,
(	2707	)	,
(	2703	)	,
(	2699	)	,
(	2695	)	,
(	2691	)	,
(	2687	)	,
(	2683	)	,
(	2679	)	,
(	2675	)	,
(	2671	)	,
(	2667	)	,
(	2663	)	,
(	2658	)	,
(	2654	)	,
(	2650	)	,
(	2646	)	,
(	2642	)	,
(	2638	)	,
(	2635	)	,
(	2631	)	,
(	2627	)	,
(	2623	)	,
(	2619	)	,
(	2615	)	,
(	2611	)	,
(	2607	)	,
(	2603	)	,
(	2599	)	,
(	2595	)	,
(	2591	)	,
(	2587	)	,
(	2583	)	,
(	2579	)	,
(	2575	)	,
(	2572	)	,
(	2568	)	,
(	2564	)	,
(	2560	)	,
(	2556	)	,
(	2552	)	,
(	2548	)	,
(	2545	)	,
(	2541	)	,
(	2537	)	,
(	2533	)	,
(	2529	)	,
(	2525	)	,
(	2522	)	,
(	2518	)	,
(	2514	)	,
(	2510	)	,
(	2506	)	,
(	2503	)	,
(	2499	)	,
(	2495	)	,
(	2491	)	,
(	2488	)	,
(	2484	)	,
(	2480	)	,
(	2476	)	,
(	2473	)	,
(	2469	)	,
(	2465	)	,
(	2461	)	,
(	2458	)	,
(	2454	)	,
(	2450	)	,
(	2446	)	,
(	2443	)	,
(	2439	)	,
(	2435	)	,
(	2432	)	,
(	2428	)	,
(	2424	)	,
(	2421	)	,
(	2417	)	,
(	2413	)	,
(	2410	)	,
(	2406	)	,
(	2403	)	,
(	2399	)	,
(	2395	)	,
(	2392	)	,
(	2388	)	,
(	2384	)	,
(	2381	)	,
(	2377	)	,
(	2374	)	,
(	2370	)	,
(	2366	)	,
(	2363	)	,
(	2359	)	,
(	2356	)	,
(	2352	)	,
(	2349	)	,
(	2345	)	,
(	2342	)	,
(	2338	)	,
(	2334	)	,
(	2331	)	,
(	2327	)	,
(	2324	)	,
(	2320	)	,
(	2317	)	,
(	2313	)	,
(	2310	)	,
(	2306	)	,
(	2303	)	,
(	2299	)	,
(	2296	)	,
(	2293	)	,
(	2289	)	,
(	2286	)	,
(	2282	)	,
(	2279	)	,
(	2275	)	,
(	2272	)	,
(	2268	)	,
(	2265	)	,
(	2262	)	,
(	2258	)	,
(	2255	)	,
(	2251	)	,
(	2248	)	,
(	2245	)	,
(	2241	)	,
(	2238	)	,
(	2234	)	,
(	2231	)	,
(	2228	)	,
(	2224	)	,
(	2221	)	,
(	2218	)	,
(	2214	)	,
(	2211	)	,
(	2208	)	,
(	2204	)	,
(	2201	)	,
(	2198	)	,
(	2194	)	,
(	2191	)	,
(	2188	)	,
(	2184	)	,
(	2181	)	,
(	2178	)	,
(	2175	)	,
(	2171	)	,
(	2168	)	,
(	2165	)	,
(	2161	)	,
(	2158	)	,
(	2155	)	,
(	2152	)	,
(	2148	)	,
(	2145	)	,
(	2142	)	,
(	2139	)	,
(	2136	)	,
(	2132	)	,
(	2129	)	,
(	2126	)	,
(	2123	)	,
(	2120	)	,
(	2116	)	,
(	2113	)	,
(	2110	)	,
(	2107	)	,
(	2104	)	,
(	2100	)	,
(	2097	)	,
(	2094	)	,
(	2091	)	,
(	2088	)	,
(	2085	)	,
(	2082	)	,
(	2078	)	,
(	2075	)	,
(	2072	)	,
(	2069	)	,
(	2066	)	,
(	2063	)	,
(	2060	)	,
(	2057	)	,
(	2054	)	,
(	2051	)	,
(	2047	)	,
(	2044	)	,
(	2041	)	,
(	2038	)	,
(	2035	)	,
(	2032	)	,
(	2029	)	,
(	2026	)	,
(	2023	)	,
(	2020	)	,
(	2017	)	,
(	2014	)	,
(	2011	)	,
(	2008	)	,
(	2005	)	,
(	2002	)	,
(	1999	)	,
(	1996	)	,
(	1993	)	,
(	1990	)	,
(	1987	)	,
(	1984	)	,
(	1981	)	,
(	1978	)	,
(	1975	)	,
(	1972	)	,
(	1969	)	,
(	1966	)	,
(	1963	)	,
(	1960	)	,
(	1957	)	,
(	1954	)	,
(	1951	)	,
(	1949	)	,
(	1946	)	,
(	1943	)	,
(	1940	)	,
(	1937	)	,
(	1934	)	,
(	1931	)	,
(	1928	)	,
(	1925	)	,
(	1922	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1900	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1886	)	,
(	1883	)	,
(	1880	)	,
(	1877	)	,
(	1874	)	,
(	1872	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1858	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1836	)	,
(	1833	)	,
(	1830	)	,
(	1827	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1809	)	,
(	1806	)	,
(	1803	)	,
(	1801	)	,
(	1798	)	,
(	1795	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1777	)	,
(	1774	)	,
(	1771	)	,
(	1769	)	,
(	1766	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1756	)	,
(	1753	)	,
(	1751	)	,
(	1748	)	,
(	1745	)	,
(	1743	)	,
(	1740	)	,
(	1738	)	,
(	1735	)	,
(	1733	)	,
(	1730	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1720	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1710	)	,
(	1707	)	,
(	1705	)	,
(	1702	)	,
(	1700	)	,
(	1697	)	,
(	1695	)	,
(	1692	)	,
(	1690	)	,
(	1687	)	,
(	1685	)	,
(	1682	)	,
(	1680	)	,
(	1678	)	,
(	1675	)	,
(	1673	)	,
(	1670	)	,
(	1668	)	,
(	1665	)	,
(	1663	)	,
(	1660	)	,
(	1658	)	,
(	1656	)	,
(	1653	)	,
(	1651	)	,
(	1648	)	,
(	1646	)	,
(	1644	)	,
(	1641	)	,
(	1639	)	,
(	1636	)	,
(	1634	)	,
(	1632	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1620	)	,
(	1617	)	,
(	1615	)	,
(	1613	)	,
(	1610	)	,
(	1608	)	,
(	1606	)	,
(	1603	)	,
(	1601	)	,
(	1599	)	,
(	1596	)	,
(	1594	)	,
(	1592	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1546	)	,
(	1544	)	,
(	1542	)	,
(	1540	)	,
(	1538	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1389	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1347	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1339	)	,
(	1338	)	,
(	1336	)	,
(	1334	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1325	)	,
(	1323	)	,
(	1321	)	,
(	1319	)	,
(	1318	)	,
(	1316	)	,
(	1314	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1303	)	,
(	1302	)	,
(	1300	)	,
(	1298	)	,
(	1296	)	,
(	1295	)	,
(	1293	)	,
(	1291	)	,
(	1289	)	,
(	1288	)	,
(	1286	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1272	)	,
(	1270	)	,
(	1269	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1257	)	,
(	1255	)	,
(	1253	)	,
(	1252	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1245	)	,
(	1244	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1235	)	,
(	1234	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1192	)	,
(	1191	)	,
(	1189	)	,
(	1188	)	,
(	1186	)	,
(	1185	)	,
(	1183	)	,
(	1182	)	,
(	1180	)	,
(	1179	)	,
(	1177	)	,
(	1175	)	,
(	1174	)	,
(	1172	)	,
(	1171	)	,
(	1169	)	,
(	1168	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1159	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1150	)	,
(	1149	)	,
(	1147	)	,
(	1146	)	,
(	1144	)	,
(	1143	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1137	)	,
(	1136	)	,
(	1134	)	,
(	1133	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1127	)	,
(	1126	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1098	)	,
(	1097	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	308	)	,
(	307	)	,
(	307	)	,
(	306	)	,
(	305	)	,
(	304	)	,
(	304	)	,
(	303	)	,
(	302	)	,
(	301	)	,
(	301	)	,
(	300	)	,
(	299	)	,
(	298	)	,
(	298	)	,
(	297	)	,
(	296	)	,
(	295	)	,
(	295	)	,
(	294	)	,
(	293	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	286	)	,
(	285	)	,
(	284	)	,
(	284	)	,
(	283	)	,
(	282	)	,
(	281	)	,
(	281	)	,
(	280	)	,
(	279	)	,
(	278	)	,
(	277	)	,
(	277	)	,
(	276	)	,
(	275	)	,
(	274	)	,
(	273	)	,
(	273	)	,
(	272	)	,
(	271	)	,
(	270	)	,
(	269	)	,
(	269	)	,
(	268	)	,
(	267	)	,
(	266	)	,
(	265	)	,
(	264	)	,
(	264	)	,
(	263	)	,
(	262	)	,
(	261	)	,
(	260	)	,
(	260	)	,
(	259	)	,
(	258	)	,
(	257	)	,
(	256	)	,
(	255	)	,
(	255	)	,
(	254	)	,
(	253	)	,
(	252	)	,
(	251	)	,
(	250	)	,
(	250	)	,
(	249	)	,
(	248	)	,
(	247	)	,
(	246	)	,
(	245	)	,
(	244	)	,
(	244	)	,
(	243	)	,
(	242	)	,
(	241	)	,
(	240	)	,
(	239	)	,
(	238	)	,
(	238	)	,
(	237	)	,
(	236	)	,
(	235	)	,
(	234	)	,
(	233	)	,
(	232	)	,
(	232	)	,
(	231	)	,
(	230	)	,
(	229	)	,
(	228	)	,
(	227	)	,
(	226	)	,
(	225	)	,
(	225	)	,
(	224	)	,
(	223	)	,
(	222	)	,
(	221	)	,
(	220	)	,
(	219	)	,
(	218	)	,
(	217	)	,
(	217	)	,
(	216	)	,
(	215	)	,
(	214	)	,
(	213	)	,
(	212	)	,
(	211	)	,
(	210	)	,
(	209	)	,
(	208	)	,
(	208	)	,
(	207	)	,
(	206	)	,
(	205	)	,
(	204	)	,
(	203	)	,
(	202	)	,
(	201	)	,
(	200	)	,
(	199	)	,
(	198	)	,
(	197	)	,
(	197	)	,
(	196	)	,
(	195	)	,
(	194	)	,
(	193	)	,
(	192	)	,
(	191	)	,
(	190	)	,
(	189	)	,
(	188	)	,
(	187	)	,
(	186	)	,
(	185	)	,
(	184	)	,
(	183	)	,
(	182	)	,
(	181	)	,
(	180	)	,
(	179	)	,
(	178	)	,
(	177	)	,
(	176	)	,
(	175	)	,
(	174	)	,
(	173	)	,
(	172	)	,
(	171	)	,
(	170	)	,
(	169	)	,
(	168	)	,
(	167	)	,
(	166	)	,
(	165	)	,
(	164	)	,
(	163	)	,
(	162	)	,
(	161	)	,
(	160	)	,
(	159	)	,
(	158	)	,
(	157	)	,
(	156	)	,
(	155	)	,
(	154	)	,
(	153	)	,
(	152	)	,
(	151	)	,
(	150	)	,
(	149	)	,
(	148	)	,
(	147	)	,
(	146	)	,
(	145	)	,
(	144	)	,
(	143	)	,
(	142	)	,
(	141	)	,
(	140	)	,
(	139	)	,
(	138	)	,
(	137	)	,
(	136	)	,
(	135	)	,
(	134	)	,
(	133	)	,
(	132	)	,
(	131	)	,
(	130	)	,
(	129	)	,
(	128	)	,
(	127	)	,
(	126	)	,
(	125	)	,
(	124	)	,
(	123	)	,
(	122	)	,
(	121	)	,
(	120	)	,
(	119	)	,
(	118	)	,
(	117	)	,
(	116	)	,
(	115	)	,
(	114	)	,
(	113	)	,
(	112	)	,
(	111	)	,
(	110	)	,
(	109	)	,
(	108	)	,
(	107	)	,
(	106	)	,
(	105	)	,
(	104	)	,
(	103	)	,
(	102	)	,
(	101	)	,
(	100	)	,
(	99	)	,
(	98	)	,
(	97	)	,
(	96	)	,
(	95	)	,
(	94	)	,
(	93	)	,
(	92	)	,
(	91	)	,
(	90	)	,
(	89	)	,
(	88	)	,
(	87	)	,
(	86	)	,
(	85	)	,
(	84	)	,
(	83	)	,
(	82	)	,
(	81	)	,
(	80	)	,
(	79	)	,
(	78	)	,
(	77	)	,
(	76	)	,
(	75	)	,
(	74	)	,
(	73	)	,
(	72	)	,
(	71	)	,
(	70	)	,
(	69	)	,
(	68	)	,
(	67	)	,
(	66	)	,
(	65	)	,
(	64	)	,
(	63	)	,
(	62	)	,
(	61	)	,
(	60	)	,
(	59	)	,
(	58	)	,
(	57	)	,
(	56	)	,
(	55	)	,
(	54	)	,
(	53	)	,
(	52	)	,
(	51	)	,
(	50	)	,
(	49	)	,
(	48	)	,
(	47	)	,
(	46	)	,
(	45	)	,
(	44	)	,
(	43	)	,
(	42	)	,
(	41	)	,
(	40	)	,
(	39	)	,
(	38	)	,
(	37	)	,
(	36	)	,
(	35	)	,
(	34	)	,
(	33	)	,
(	32	)	,
(	31	)	,
(	30	)	,
(	29	)	,
(	28	)	,
(	27	)	,
(	26	)	,
(	25	)	,
(	24	)	,
(	23	)	,
(	22	)	,
(	21	)	,
(	20	)	,
(	19	)	,
(	18	)	,
(	17	)	,
(	16	)	,
(	15	)	,
(	14	)	,
(	13	)	,
(	12	)	,
(	11	)	,
(	10	)	,
(	9	)	,
(	8	)	,
(	7	)	,
(	6	)	,
(	5	)	,
(	4	)	,
(	3	)	,
(	2	)	,
(	1	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	




);


end package LUT_pkg;
