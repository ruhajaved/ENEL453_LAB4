library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LED_Flash_LUT_pkg is
 
 type my_array is array (4095 downto 0) of integer;
 constant DtoP_LUT : my_array := (
 
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	60000	)	,
(	59985	)	,
(	59970	)	,
(	59955	)	,
(	59940	)	,
(	59925	)	,
(	59910	)	,
(	59895	)	,
(	59880	)	,
(	59865	)	,
(	59850	)	,
(	59835	)	,
(	59820	)	,
(	59805	)	,
(	59790	)	,
(	59775	)	,
(	59760	)	,
(	59745	)	,
(	59730	)	,
(	59715	)	,
(	59700	)	,
(	59685	)	,
(	59670	)	,
(	59655	)	,
(	59640	)	,
(	59625	)	,
(	59610	)	,
(	59595	)	,
(	59580	)	,
(	59565	)	,
(	59550	)	,
(	59535	)	,
(	59520	)	,
(	59505	)	,
(	59490	)	,
(	59475	)	,
(	59460	)	,
(	59445	)	,
(	59430	)	,
(	59415	)	,
(	59400	)	,
(	59385	)	,
(	59370	)	,
(	59355	)	,
(	59340	)	,
(	59325	)	,
(	59310	)	,
(	59295	)	,
(	59280	)	,
(	59265	)	,
(	59250	)	,
(	59235	)	,
(	59220	)	,
(	59205	)	,
(	59190	)	,
(	59175	)	,
(	59160	)	,
(	59145	)	,
(	59130	)	,
(	59115	)	,
(	59100	)	,
(	59085	)	,
(	59070	)	,
(	59055	)	,
(	59040	)	,
(	59025	)	,
(	59010	)	,
(	58995	)	,
(	58980	)	,
(	58965	)	,
(	58950	)	,
(	58935	)	,
(	58920	)	,
(	58905	)	,
(	58890	)	,
(	58875	)	,
(	58860	)	,
(	58845	)	,
(	58830	)	,
(	58815	)	,
(	58800	)	,
(	58785	)	,
(	58770	)	,
(	58755	)	,
(	58740	)	,
(	58725	)	,
(	58710	)	,
(	58695	)	,
(	58680	)	,
(	58665	)	,
(	58650	)	,
(	58635	)	,
(	58620	)	,
(	58605	)	,
(	58590	)	,
(	58575	)	,
(	58560	)	,
(	58545	)	,
(	58530	)	,
(	58515	)	,
(	58500	)	,
(	58485	)	,
(	58470	)	,
(	58455	)	,
(	58440	)	,
(	58425	)	,
(	58410	)	,
(	58395	)	,
(	58380	)	,
(	58365	)	,
(	58350	)	,
(	58335	)	,
(	58320	)	,
(	58305	)	,
(	58290	)	,
(	58275	)	,
(	58260	)	,
(	58245	)	,
(	58230	)	,
(	58215	)	,
(	58200	)	,
(	58185	)	,
(	58170	)	,
(	58155	)	,
(	58140	)	,
(	58125	)	,
(	58110	)	,
(	58095	)	,
(	58080	)	,
(	58065	)	,
(	58050	)	,
(	58035	)	,
(	58020	)	,
(	58005	)	,
(	57990	)	,
(	57975	)	,
(	57960	)	,
(	57945	)	,
(	57930	)	,
(	57915	)	,
(	57900	)	,
(	57885	)	,
(	57870	)	,
(	57855	)	,
(	57840	)	,
(	57825	)	,
(	57810	)	,
(	57795	)	,
(	57780	)	,
(	57765	)	,
(	57750	)	,
(	57735	)	,
(	57720	)	,
(	57705	)	,
(	57690	)	,
(	57675	)	,
(	57660	)	,
(	57645	)	,
(	57630	)	,
(	57615	)	,
(	57600	)	,
(	57585	)	,
(	57570	)	,
(	57555	)	,
(	57540	)	,
(	57525	)	,
(	57510	)	,
(	57495	)	,
(	57480	)	,
(	57465	)	,
(	57450	)	,
(	57435	)	,
(	57420	)	,
(	57405	)	,
(	57390	)	,
(	57375	)	,
(	57360	)	,
(	57345	)	,
(	57330	)	,
(	57315	)	,
(	57300	)	,
(	57285	)	,
(	57270	)	,
(	57255	)	,
(	57240	)	,
(	57225	)	,
(	57210	)	,
(	57195	)	,
(	57180	)	,
(	57165	)	,
(	57150	)	,
(	57135	)	,
(	57120	)	,
(	57105	)	,
(	57090	)	,
(	57075	)	,
(	57060	)	,
(	57045	)	,
(	57030	)	,
(	57015	)	,
(	57000	)	,
(	56985	)	,
(	56970	)	,
(	56955	)	,
(	56940	)	,
(	56925	)	,
(	56910	)	,
(	56895	)	,
(	56880	)	,
(	56865	)	,
(	56850	)	,
(	56835	)	,
(	56820	)	,
(	56805	)	,
(	56790	)	,
(	56775	)	,
(	56760	)	,
(	56745	)	,
(	56730	)	,
(	56715	)	,
(	56700	)	,
(	56685	)	,
(	56670	)	,
(	56655	)	,
(	56640	)	,
(	56625	)	,
(	56610	)	,
(	56595	)	,
(	56580	)	,
(	56565	)	,
(	56550	)	,
(	56535	)	,
(	56520	)	,
(	56505	)	,
(	56490	)	,
(	56475	)	,
(	56460	)	,
(	56445	)	,
(	56430	)	,
(	56415	)	,
(	56400	)	,
(	56385	)	,
(	56370	)	,
(	56355	)	,
(	56340	)	,
(	56325	)	,
(	56310	)	,
(	56295	)	,
(	56280	)	,
(	56265	)	,
(	56250	)	,
(	56235	)	,
(	56220	)	,
(	56205	)	,
(	56190	)	,
(	56175	)	,
(	56160	)	,
(	56145	)	,
(	56130	)	,
(	56115	)	,
(	56100	)	,
(	56085	)	,
(	56070	)	,
(	56055	)	,
(	56040	)	,
(	56025	)	,
(	56010	)	,
(	55995	)	,
(	55980	)	,
(	55965	)	,
(	55950	)	,
(	55935	)	,
(	55920	)	,
(	55905	)	,
(	55890	)	,
(	55875	)	,
(	55860	)	,
(	55845	)	,
(	55830	)	,
(	55815	)	,
(	55800	)	,
(	55785	)	,
(	55770	)	,
(	55755	)	,
(	55740	)	,
(	55725	)	,
(	55710	)	,
(	55695	)	,
(	55680	)	,
(	55665	)	,
(	55650	)	,
(	55635	)	,
(	55620	)	,
(	55605	)	,
(	55590	)	,
(	55575	)	,
(	55560	)	,
(	55545	)	,
(	55530	)	,
(	55515	)	,
(	55500	)	,
(	55485	)	,
(	55470	)	,
(	55455	)	,
(	55440	)	,
(	55425	)	,
(	55410	)	,
(	55395	)	,
(	55380	)	,
(	55365	)	,
(	55350	)	,
(	55335	)	,
(	55320	)	,
(	55305	)	,
(	55290	)	,
(	55275	)	,
(	55260	)	,
(	55245	)	,
(	55230	)	,
(	55215	)	,
(	55200	)	,
(	55185	)	,
(	55170	)	,
(	55155	)	,
(	55140	)	,
(	55125	)	,
(	55110	)	,
(	55095	)	,
(	55080	)	,
(	55065	)	,
(	55050	)	,
(	55035	)	,
(	55020	)	,
(	55005	)	,
(	54990	)	,
(	54975	)	,
(	54960	)	,
(	54945	)	,
(	54930	)	,
(	54915	)	,
(	54900	)	,
(	54885	)	,
(	54870	)	,
(	54855	)	,
(	54840	)	,
(	54825	)	,
(	54810	)	,
(	54795	)	,
(	54780	)	,
(	54765	)	,
(	54750	)	,
(	54735	)	,
(	54720	)	,
(	54705	)	,
(	54690	)	,
(	54675	)	,
(	54660	)	,
(	54645	)	,
(	54630	)	,
(	54615	)	,
(	54600	)	,
(	54585	)	,
(	54570	)	,
(	54555	)	,
(	54540	)	,
(	54525	)	,
(	54510	)	,
(	54495	)	,
(	54480	)	,
(	54465	)	,
(	54450	)	,
(	54435	)	,
(	54420	)	,
(	54405	)	,
(	54390	)	,
(	54375	)	,
(	54360	)	,
(	54345	)	,
(	54330	)	,
(	54315	)	,
(	54300	)	,
(	54285	)	,
(	54270	)	,
(	54255	)	,
(	54240	)	,
(	54225	)	,
(	54210	)	,
(	54195	)	,
(	54180	)	,
(	54165	)	,
(	54150	)	,
(	54135	)	,
(	54120	)	,
(	54105	)	,
(	54090	)	,
(	54075	)	,
(	54060	)	,
(	54045	)	,
(	54030	)	,
(	54015	)	,
(	54000	)	,
(	53985	)	,
(	53970	)	,
(	53955	)	,
(	53940	)	,
(	53925	)	,
(	53910	)	,
(	53895	)	,
(	53880	)	,
(	53865	)	,
(	53850	)	,
(	53835	)	,
(	53820	)	,
(	53805	)	,
(	53790	)	,
(	53775	)	,
(	53760	)	,
(	53745	)	,
(	53730	)	,
(	53715	)	,
(	53700	)	,
(	53685	)	,
(	53670	)	,
(	53655	)	,
(	53640	)	,
(	53625	)	,
(	53610	)	,
(	53595	)	,
(	53580	)	,
(	53565	)	,
(	53550	)	,
(	53535	)	,
(	53520	)	,
(	53505	)	,
(	53490	)	,
(	53475	)	,
(	53460	)	,
(	53445	)	,
(	53430	)	,
(	53415	)	,
(	53400	)	,
(	53385	)	,
(	53370	)	,
(	53355	)	,
(	53340	)	,
(	53325	)	,
(	53310	)	,
(	53295	)	,
(	53280	)	,
(	53265	)	,
(	53250	)	,
(	53235	)	,
(	53220	)	,
(	53205	)	,
(	53190	)	,
(	53175	)	,
(	53160	)	,
(	53145	)	,
(	53130	)	,
(	53115	)	,
(	53100	)	,
(	53085	)	,
(	53070	)	,
(	53055	)	,
(	53040	)	,
(	53025	)	,
(	53010	)	,
(	52995	)	,
(	52980	)	,
(	52965	)	,
(	52950	)	,
(	52935	)	,
(	52920	)	,
(	52905	)	,
(	52890	)	,
(	52875	)	,
(	52860	)	,
(	52845	)	,
(	52830	)	,
(	52815	)	,
(	52800	)	,
(	52785	)	,
(	52770	)	,
(	52755	)	,
(	52740	)	,
(	52725	)	,
(	52710	)	,
(	52695	)	,
(	52680	)	,
(	52665	)	,
(	52650	)	,
(	52635	)	,
(	52620	)	,
(	52605	)	,
(	52590	)	,
(	52575	)	,
(	52560	)	,
(	52545	)	,
(	52530	)	,
(	52515	)	,
(	52500	)	,
(	52485	)	,
(	52470	)	,
(	52455	)	,
(	52440	)	,
(	52425	)	,
(	52410	)	,
(	52395	)	,
(	52380	)	,
(	52365	)	,
(	52350	)	,
(	52335	)	,
(	52320	)	,
(	52305	)	,
(	52290	)	,
(	52275	)	,
(	52260	)	,
(	52245	)	,
(	52230	)	,
(	52215	)	,
(	52200	)	,
(	52185	)	,
(	52170	)	,
(	52155	)	,
(	52140	)	,
(	52125	)	,
(	52110	)	,
(	52095	)	,
(	52080	)	,
(	52065	)	,
(	52050	)	,
(	52035	)	,
(	52020	)	,
(	52005	)	,
(	51990	)	,
(	51975	)	,
(	51960	)	,
(	51945	)	,
(	51930	)	,
(	51915	)	,
(	51900	)	,
(	51885	)	,
(	51870	)	,
(	51855	)	,
(	51840	)	,
(	51825	)	,
(	51810	)	,
(	51795	)	,
(	51780	)	,
(	51765	)	,
(	51750	)	,
(	51735	)	,
(	51720	)	,
(	51705	)	,
(	51690	)	,
(	51675	)	,
(	51660	)	,
(	51645	)	,
(	51630	)	,
(	51615	)	,
(	51600	)	,
(	51585	)	,
(	51570	)	,
(	51555	)	,
(	51540	)	,
(	51525	)	,
(	51510	)	,
(	51495	)	,
(	51480	)	,
(	51465	)	,
(	51450	)	,
(	51435	)	,
(	51420	)	,
(	51405	)	,
(	51390	)	,
(	51375	)	,
(	51360	)	,
(	51345	)	,
(	51330	)	,
(	51315	)	,
(	51300	)	,
(	51285	)	,
(	51270	)	,
(	51255	)	,
(	51240	)	,
(	51225	)	,
(	51210	)	,
(	51195	)	,
(	51180	)	,
(	51165	)	,
(	51150	)	,
(	51135	)	,
(	51120	)	,
(	51105	)	,
(	51090	)	,
(	51075	)	,
(	51060	)	,
(	51045	)	,
(	51030	)	,
(	51015	)	,
(	51000	)	,
(	50985	)	,
(	50970	)	,
(	50955	)	,
(	50940	)	,
(	50925	)	,
(	50910	)	,
(	50895	)	,
(	50880	)	,
(	50865	)	,
(	50850	)	,
(	50835	)	,
(	50820	)	,
(	50805	)	,
(	50790	)	,
(	50775	)	,
(	50760	)	,
(	50745	)	,
(	50730	)	,
(	50715	)	,
(	50700	)	,
(	50685	)	,
(	50670	)	,
(	50655	)	,
(	50640	)	,
(	50625	)	,
(	50610	)	,
(	50595	)	,
(	50580	)	,
(	50565	)	,
(	50550	)	,
(	50535	)	,
(	50520	)	,
(	50505	)	,
(	50490	)	,
(	50475	)	,
(	50460	)	,
(	50445	)	,
(	50430	)	,
(	50415	)	,
(	50400	)	,
(	50385	)	,
(	50370	)	,
(	50355	)	,
(	50340	)	,
(	50325	)	,
(	50310	)	,
(	50295	)	,
(	50280	)	,
(	50265	)	,
(	50250	)	,
(	50235	)	,
(	50220	)	,
(	50205	)	,
(	50190	)	,
(	50175	)	,
(	50160	)	,
(	50145	)	,
(	50130	)	,
(	50115	)	,
(	50100	)	,
(	50085	)	,
(	50070	)	,
(	50055	)	,
(	50040	)	,
(	50025	)	,
(	50010	)	,
(	49995	)	,
(	49980	)	,
(	49965	)	,
(	49950	)	,
(	49935	)	,
(	49920	)	,
(	49905	)	,
(	49890	)	,
(	49875	)	,
(	49860	)	,
(	49845	)	,
(	49830	)	,
(	49815	)	,
(	49800	)	,
(	49785	)	,
(	49770	)	,
(	49755	)	,
(	49740	)	,
(	49725	)	,
(	49710	)	,
(	49695	)	,
(	49680	)	,
(	49665	)	,
(	49650	)	,
(	49635	)	,
(	49620	)	,
(	49605	)	,
(	49590	)	,
(	49575	)	,
(	49560	)	,
(	49545	)	,
(	49530	)	,
(	49515	)	,
(	49500	)	,
(	49485	)	,
(	49470	)	,
(	49455	)	,
(	49440	)	,
(	49425	)	,
(	49410	)	,
(	49395	)	,
(	49380	)	,
(	49365	)	,
(	49350	)	,
(	49335	)	,
(	49320	)	,
(	49305	)	,
(	49290	)	,
(	49275	)	,
(	49260	)	,
(	49245	)	,
(	49230	)	,
(	49215	)	,
(	49200	)	,
(	49185	)	,
(	49170	)	,
(	49155	)	,
(	49140	)	,
(	49125	)	,
(	49110	)	,
(	49095	)	,
(	49080	)	,
(	49065	)	,
(	49050	)	,
(	49035	)	,
(	49020	)	,
(	49005	)	,
(	48990	)	,
(	48975	)	,
(	48960	)	,
(	48945	)	,
(	48930	)	,
(	48915	)	,
(	48900	)	,
(	48885	)	,
(	48870	)	,
(	48855	)	,
(	48840	)	,
(	48825	)	,
(	48810	)	,
(	48795	)	,
(	48780	)	,
(	48765	)	,
(	48750	)	,
(	48735	)	,
(	48720	)	,
(	48705	)	,
(	48690	)	,
(	48675	)	,
(	48660	)	,
(	48645	)	,
(	48630	)	,
(	48615	)	,
(	48600	)	,
(	48585	)	,
(	48570	)	,
(	48555	)	,
(	48540	)	,
(	48525	)	,
(	48510	)	,
(	48495	)	,
(	48480	)	,
(	48465	)	,
(	48450	)	,
(	48435	)	,
(	48420	)	,
(	48405	)	,
(	48390	)	,
(	48375	)	,
(	48360	)	,
(	48345	)	,
(	48330	)	,
(	48315	)	,
(	48300	)	,
(	48285	)	,
(	48270	)	,
(	48255	)	,
(	48240	)	,
(	48225	)	,
(	48210	)	,
(	48195	)	,
(	48180	)	,
(	48165	)	,
(	48150	)	,
(	48135	)	,
(	48120	)	,
(	48105	)	,
(	48090	)	,
(	48075	)	,
(	48060	)	,
(	48045	)	,
(	48030	)	,
(	48015	)	,
(	48000	)	,
(	47985	)	,
(	47970	)	,
(	47955	)	,
(	47940	)	,
(	47925	)	,
(	47910	)	,
(	47895	)	,
(	47880	)	,
(	47865	)	,
(	47850	)	,
(	47835	)	,
(	47820	)	,
(	47805	)	,
(	47790	)	,
(	47775	)	,
(	47760	)	,
(	47745	)	,
(	47730	)	,
(	47715	)	,
(	47700	)	,
(	47685	)	,
(	47670	)	,
(	47655	)	,
(	47640	)	,
(	47625	)	,
(	47610	)	,
(	47595	)	,
(	47580	)	,
(	47565	)	,
(	47550	)	,
(	47535	)	,
(	47520	)	,
(	47505	)	,
(	47490	)	,
(	47475	)	,
(	47460	)	,
(	47445	)	,
(	47430	)	,
(	47415	)	,
(	47400	)	,
(	47385	)	,
(	47370	)	,
(	47355	)	,
(	47340	)	,
(	47325	)	,
(	47310	)	,
(	47295	)	,
(	47280	)	,
(	47265	)	,
(	47250	)	,
(	47235	)	,
(	47220	)	,
(	47205	)	,
(	47190	)	,
(	47175	)	,
(	47160	)	,
(	47145	)	,
(	47130	)	,
(	47115	)	,
(	47100	)	,
(	47085	)	,
(	47070	)	,
(	47055	)	,
(	47040	)	,
(	47025	)	,
(	47010	)	,
(	46995	)	,
(	46980	)	,
(	46965	)	,
(	46950	)	,
(	46935	)	,
(	46920	)	,
(	46905	)	,
(	46890	)	,
(	46875	)	,
(	46860	)	,
(	46845	)	,
(	46830	)	,
(	46815	)	,
(	46800	)	,
(	46785	)	,
(	46770	)	,
(	46755	)	,
(	46740	)	,
(	46725	)	,
(	46710	)	,
(	46695	)	,
(	46680	)	,
(	46665	)	,
(	46650	)	,
(	46635	)	,
(	46620	)	,
(	46605	)	,
(	46590	)	,
(	46575	)	,
(	46560	)	,
(	46545	)	,
(	46530	)	,
(	46515	)	,
(	46500	)	,
(	46485	)	,
(	46470	)	,
(	46455	)	,
(	46440	)	,
(	46425	)	,
(	46410	)	,
(	46395	)	,
(	46380	)	,
(	46365	)	,
(	46350	)	,
(	46335	)	,
(	46320	)	,
(	46305	)	,
(	46290	)	,
(	46275	)	,
(	46260	)	,
(	46245	)	,
(	46230	)	,
(	46215	)	,
(	46200	)	,
(	46185	)	,
(	46170	)	,
(	46155	)	,
(	46140	)	,
(	46125	)	,
(	46110	)	,
(	46095	)	,
(	46080	)	,
(	46065	)	,
(	46050	)	,
(	46035	)	,
(	46020	)	,
(	46005	)	,
(	45990	)	,
(	45975	)	,
(	45960	)	,
(	45945	)	,
(	45930	)	,
(	45915	)	,
(	45900	)	,
(	45885	)	,
(	45870	)	,
(	45855	)	,
(	45840	)	,
(	45825	)	,
(	45810	)	,
(	45795	)	,
(	45780	)	,
(	45765	)	,
(	45750	)	,
(	45735	)	,
(	45720	)	,
(	45705	)	,
(	45690	)	,
(	45675	)	,
(	45660	)	,
(	45645	)	,
(	45630	)	,
(	45615	)	,
(	45600	)	,
(	45585	)	,
(	45570	)	,
(	45555	)	,
(	45540	)	,
(	45525	)	,
(	45510	)	,
(	45495	)	,
(	45480	)	,
(	45465	)	,
(	45450	)	,
(	45435	)	,
(	45420	)	,
(	45405	)	,
(	45390	)	,
(	45375	)	,
(	45360	)	,
(	45345	)	,
(	45330	)	,
(	45315	)	,
(	45300	)	,
(	45285	)	,
(	45270	)	,
(	45255	)	,
(	45240	)	,
(	45225	)	,
(	45210	)	,
(	45195	)	,
(	45180	)	,
(	45165	)	,
(	45150	)	,
(	45135	)	,
(	45120	)	,
(	45105	)	,
(	45090	)	,
(	45075	)	,
(	45060	)	,
(	45045	)	,
(	45030	)	,
(	45015	)	,
(	45000	)	,
(	44985	)	,
(	44970	)	,
(	44955	)	,
(	44940	)	,
(	44925	)	,
(	44910	)	,
(	44895	)	,
(	44880	)	,
(	44865	)	,
(	44850	)	,
(	44835	)	,
(	44820	)	,
(	44805	)	,
(	44790	)	,
(	44775	)	,
(	44760	)	,
(	44745	)	,
(	44730	)	,
(	44715	)	,
(	44700	)	,
(	44685	)	,
(	44670	)	,
(	44655	)	,
(	44640	)	,
(	44625	)	,
(	44610	)	,
(	44595	)	,
(	44580	)	,
(	44565	)	,
(	44550	)	,
(	44535	)	,
(	44520	)	,
(	44505	)	,
(	44490	)	,
(	44475	)	,
(	44460	)	,
(	44445	)	,
(	44430	)	,
(	44415	)	,
(	44400	)	,
(	44385	)	,
(	44370	)	,
(	44355	)	,
(	44340	)	,
(	44325	)	,
(	44310	)	,
(	44295	)	,
(	44280	)	,
(	44265	)	,
(	44250	)	,
(	44235	)	,
(	44220	)	,
(	44205	)	,
(	44190	)	,
(	44175	)	,
(	44160	)	,
(	44145	)	,
(	44130	)	,
(	44115	)	,
(	44100	)	,
(	44085	)	,
(	44070	)	,
(	44055	)	,
(	44040	)	,
(	44025	)	,
(	44010	)	,
(	43995	)	,
(	43980	)	,
(	43965	)	,
(	43950	)	,
(	43935	)	,
(	43920	)	,
(	43905	)	,
(	43890	)	,
(	43875	)	,
(	43860	)	,
(	43845	)	,
(	43830	)	,
(	43815	)	,
(	43800	)	,
(	43785	)	,
(	43770	)	,
(	43755	)	,
(	43740	)	,
(	43725	)	,
(	43710	)	,
(	43695	)	,
(	43680	)	,
(	43665	)	,
(	43650	)	,
(	43635	)	,
(	43620	)	,
(	43605	)	,
(	43590	)	,
(	43575	)	,
(	43560	)	,
(	43545	)	,
(	43530	)	,
(	43515	)	,
(	43500	)	,
(	43485	)	,
(	43470	)	,
(	43455	)	,
(	43440	)	,
(	43425	)	,
(	43410	)	,
(	43395	)	,
(	43380	)	,
(	43365	)	,
(	43350	)	,
(	43335	)	,
(	43320	)	,
(	43305	)	,
(	43290	)	,
(	43275	)	,
(	43260	)	,
(	43245	)	,
(	43230	)	,
(	43215	)	,
(	43200	)	,
(	43185	)	,
(	43170	)	,
(	43155	)	,
(	43140	)	,
(	43125	)	,
(	43110	)	,
(	43095	)	,
(	43080	)	,
(	43065	)	,
(	43050	)	,
(	43035	)	,
(	43020	)	,
(	43005	)	,
(	42990	)	,
(	42975	)	,
(	42960	)	,
(	42945	)	,
(	42930	)	,
(	42915	)	,
(	42900	)	,
(	42885	)	,
(	42870	)	,
(	42855	)	,
(	42840	)	,
(	42825	)	,
(	42810	)	,
(	42795	)	,
(	42780	)	,
(	42765	)	,
(	42750	)	,
(	42735	)	,
(	42720	)	,
(	42705	)	,
(	42690	)	,
(	42675	)	,
(	42660	)	,
(	42645	)	,
(	42630	)	,
(	42615	)	,
(	42600	)	,
(	42585	)	,
(	42570	)	,
(	42555	)	,
(	42540	)	,
(	42525	)	,
(	42510	)	,
(	42495	)	,
(	42480	)	,
(	42465	)	,
(	42450	)	,
(	42435	)	,
(	42420	)	,
(	42405	)	,
(	42390	)	,
(	42375	)	,
(	42360	)	,
(	42345	)	,
(	42330	)	,
(	42315	)	,
(	42300	)	,
(	42285	)	,
(	42270	)	,
(	42255	)	,
(	42240	)	,
(	42225	)	,
(	42210	)	,
(	42195	)	,
(	42180	)	,
(	42165	)	,
(	42150	)	,
(	42135	)	,
(	42120	)	,
(	42105	)	,
(	42090	)	,
(	42075	)	,
(	42060	)	,
(	42045	)	,
(	42030	)	,
(	42015	)	,
(	42000	)	,
(	41985	)	,
(	41970	)	,
(	41955	)	,
(	41940	)	,
(	41925	)	,
(	41910	)	,
(	41895	)	,
(	41880	)	,
(	41865	)	,
(	41850	)	,
(	41835	)	,
(	41820	)	,
(	41805	)	,
(	41790	)	,
(	41775	)	,
(	41760	)	,
(	41745	)	,
(	41730	)	,
(	41715	)	,
(	41700	)	,
(	41685	)	,
(	41670	)	,
(	41655	)	,
(	41640	)	,
(	41625	)	,
(	41610	)	,
(	41595	)	,
(	41580	)	,
(	41565	)	,
(	41550	)	,
(	41535	)	,
(	41520	)	,
(	41505	)	,
(	41490	)	,
(	41475	)	,
(	41460	)	,
(	41445	)	,
(	41430	)	,
(	41415	)	,
(	41400	)	,
(	41385	)	,
(	41370	)	,
(	41355	)	,
(	41340	)	,
(	41325	)	,
(	41310	)	,
(	41295	)	,
(	41280	)	,
(	41265	)	,
(	41250	)	,
(	41235	)	,
(	41220	)	,
(	41205	)	,
(	41190	)	,
(	41175	)	,
(	41160	)	,
(	41145	)	,
(	41130	)	,
(	41115	)	,
(	41100	)	,
(	41085	)	,
(	41070	)	,
(	41055	)	,
(	41040	)	,
(	41025	)	,
(	41010	)	,
(	40995	)	,
(	40980	)	,
(	40965	)	,
(	40950	)	,
(	40935	)	,
(	40920	)	,
(	40905	)	,
(	40890	)	,
(	40875	)	,
(	40860	)	,
(	40845	)	,
(	40830	)	,
(	40815	)	,
(	40800	)	,
(	40785	)	,
(	40770	)	,
(	40755	)	,
(	40740	)	,
(	40725	)	,
(	40710	)	,
(	40695	)	,
(	40680	)	,
(	40665	)	,
(	40650	)	,
(	40635	)	,
(	40620	)	,
(	40605	)	,
(	40590	)	,
(	40575	)	,
(	40560	)	,
(	40545	)	,
(	40530	)	,
(	40515	)	,
(	40500	)	,
(	40485	)	,
(	40470	)	,
(	40455	)	,
(	40440	)	,
(	40425	)	,
(	40410	)	,
(	40395	)	,
(	40380	)	,
(	40365	)	,
(	40350	)	,
(	40335	)	,
(	40320	)	,
(	40305	)	,
(	40290	)	,
(	40275	)	,
(	40260	)	,
(	40245	)	,
(	40230	)	,
(	40215	)	,
(	40200	)	,
(	40185	)	,
(	40170	)	,
(	40155	)	,
(	40140	)	,
(	40125	)	,
(	40110	)	,
(	40095	)	,
(	40080	)	,
(	40065	)	,
(	40050	)	,
(	40035	)	,
(	40020	)	,
(	40005	)	,
(	39990	)	,
(	39975	)	,
(	39960	)	,
(	39945	)	,
(	39930	)	,
(	39915	)	,
(	39900	)	,
(	39885	)	,
(	39870	)	,
(	39855	)	,
(	39840	)	,
(	39825	)	,
(	39810	)	,
(	39795	)	,
(	39780	)	,
(	39765	)	,
(	39750	)	,
(	39735	)	,
(	39720	)	,
(	39705	)	,
(	39690	)	,
(	39675	)	,
(	39660	)	,
(	39645	)	,
(	39630	)	,
(	39615	)	,
(	39600	)	,
(	39585	)	,
(	39570	)	,
(	39555	)	,
(	39540	)	,
(	39525	)	,
(	39510	)	,
(	39495	)	,
(	39480	)	,
(	39465	)	,
(	39450	)	,
(	39435	)	,
(	39420	)	,
(	39405	)	,
(	39390	)	,
(	39375	)	,
(	39360	)	,
(	39345	)	,
(	39330	)	,
(	39315	)	,
(	39300	)	,
(	39285	)	,
(	39270	)	,
(	39255	)	,
(	39240	)	,
(	39225	)	,
(	39210	)	,
(	39195	)	,
(	39180	)	,
(	39165	)	,
(	39150	)	,
(	39135	)	,
(	39120	)	,
(	39105	)	,
(	39090	)	,
(	39075	)	,
(	39060	)	,
(	39045	)	,
(	39030	)	,
(	39015	)	,
(	39000	)	,
(	38985	)	,
(	38970	)	,
(	38955	)	,
(	38940	)	,
(	38925	)	,
(	38910	)	,
(	38895	)	,
(	38880	)	,
(	38865	)	,
(	38850	)	,
(	38835	)	,
(	38820	)	,
(	38805	)	,
(	38790	)	,
(	38775	)	,
(	38760	)	,
(	38745	)	,
(	38730	)	,
(	38715	)	,
(	38700	)	,
(	38685	)	,
(	38670	)	,
(	38655	)	,
(	38640	)	,
(	38625	)	,
(	38610	)	,
(	38595	)	,
(	38580	)	,
(	38565	)	,
(	38550	)	,
(	38535	)	,
(	38520	)	,
(	38505	)	,
(	38490	)	,
(	38475	)	,
(	38460	)	,
(	38445	)	,
(	38430	)	,
(	38415	)	,
(	38400	)	,
(	38385	)	,
(	38370	)	,
(	38355	)	,
(	38340	)	,
(	38325	)	,
(	38310	)	,
(	38295	)	,
(	38280	)	,
(	38265	)	,
(	38250	)	,
(	38235	)	,
(	38220	)	,
(	38205	)	,
(	38190	)	,
(	38175	)	,
(	38160	)	,
(	38145	)	,
(	38130	)	,
(	38115	)	,
(	38100	)	,
(	38085	)	,
(	38070	)	,
(	38055	)	,
(	38040	)	,
(	38025	)	,
(	38010	)	,
(	37995	)	,
(	37980	)	,
(	37965	)	,
(	37950	)	,
(	37935	)	,
(	37920	)	,
(	37905	)	,
(	37890	)	,
(	37875	)	,
(	37860	)	,
(	37845	)	,
(	37830	)	,
(	37815	)	,
(	37800	)	,
(	37785	)	,
(	37770	)	,
(	37755	)	,
(	37740	)	,
(	37725	)	,
(	37710	)	,
(	37695	)	,
(	37680	)	,
(	37665	)	,
(	37650	)	,
(	37635	)	,
(	37620	)	,
(	37605	)	,
(	37590	)	,
(	37575	)	,
(	37560	)	,
(	37545	)	,
(	37530	)	,
(	37515	)	,
(	37500	)	,
(	37485	)	,
(	37470	)	,
(	37455	)	,
(	37440	)	,
(	37425	)	,
(	37410	)	,
(	37395	)	,
(	37380	)	,
(	37365	)	,
(	37350	)	,
(	37335	)	,
(	37320	)	,
(	37305	)	,
(	37290	)	,
(	37275	)	,
(	37260	)	,
(	37245	)	,
(	37230	)	,
(	37215	)	,
(	37200	)	,
(	37185	)	,
(	37170	)	,
(	37155	)	,
(	37140	)	,
(	37125	)	,
(	37110	)	,
(	37095	)	,
(	37080	)	,
(	37065	)	,
(	37050	)	,
(	37035	)	,
(	37020	)	,
(	37005	)	,
(	36990	)	,
(	36975	)	,
(	36960	)	,
(	36945	)	,
(	36930	)	,
(	36915	)	,
(	36900	)	,
(	36885	)	,
(	36870	)	,
(	36855	)	,
(	36840	)	,
(	36825	)	,
(	36810	)	,
(	36795	)	,
(	36780	)	,
(	36765	)	,
(	36750	)	,
(	36735	)	,
(	36720	)	,
(	36705	)	,
(	36690	)	,
(	36675	)	,
(	36660	)	,
(	36645	)	,
(	36630	)	,
(	36615	)	,
(	36600	)	,
(	36585	)	,
(	36570	)	,
(	36555	)	,
(	36540	)	,
(	36525	)	,
(	36510	)	,
(	36495	)	,
(	36480	)	,
(	36465	)	,
(	36450	)	,
(	36435	)	,
(	36420	)	,
(	36405	)	,
(	36390	)	,
(	36375	)	,
(	36360	)	,
(	36345	)	,
(	36330	)	,
(	36315	)	,
(	36300	)	,
(	36285	)	,
(	36270	)	,
(	36255	)	,
(	36240	)	,
(	36225	)	,
(	36210	)	,
(	36195	)	,
(	36180	)	,
(	36165	)	,
(	36150	)	,
(	36135	)	,
(	36120	)	,
(	36105	)	,
(	36090	)	,
(	36075	)	,
(	36060	)	,
(	36045	)	,
(	36030	)	,
(	36015	)	,
(	36000	)	,
(	35985	)	,
(	35970	)	,
(	35955	)	,
(	35940	)	,
(	35925	)	,
(	35910	)	,
(	35895	)	,
(	35880	)	,
(	35865	)	,
(	35850	)	,
(	35835	)	,
(	35820	)	,
(	35805	)	,
(	35790	)	,
(	35775	)	,
(	35760	)	,
(	35745	)	,
(	35730	)	,
(	35715	)	,
(	35700	)	,
(	35685	)	,
(	35670	)	,
(	35655	)	,
(	35640	)	,
(	35625	)	,
(	35610	)	,
(	35595	)	,
(	35580	)	,
(	35565	)	,
(	35550	)	,
(	35535	)	,
(	35520	)	,
(	35505	)	,
(	35490	)	,
(	35475	)	,
(	35460	)	,
(	35445	)	,
(	35430	)	,
(	35415	)	,
(	35400	)	,
(	35385	)	,
(	35370	)	,
(	35355	)	,
(	35340	)	,
(	35325	)	,
(	35310	)	,
(	35295	)	,
(	35280	)	,
(	35265	)	,
(	35250	)	,
(	35235	)	,
(	35220	)	,
(	35205	)	,
(	35190	)	,
(	35175	)	,
(	35160	)	,
(	35145	)	,
(	35130	)	,
(	35115	)	,
(	35100	)	,
(	35085	)	,
(	35070	)	,
(	35055	)	,
(	35040	)	,
(	35025	)	,
(	35010	)	,
(	34995	)	,
(	34980	)	,
(	34965	)	,
(	34950	)	,
(	34935	)	,
(	34920	)	,
(	34905	)	,
(	34890	)	,
(	34875	)	,
(	34860	)	,
(	34845	)	,
(	34830	)	,
(	34815	)	,
(	34800	)	,
(	34785	)	,
(	34770	)	,
(	34755	)	,
(	34740	)	,
(	34725	)	,
(	34710	)	,
(	34695	)	,
(	34680	)	,
(	34665	)	,
(	34650	)	,
(	34635	)	,
(	34620	)	,
(	34605	)	,
(	34590	)	,
(	34575	)	,
(	34560	)	,
(	34545	)	,
(	34530	)	,
(	34515	)	,
(	34500	)	,
(	34485	)	,
(	34470	)	,
(	34455	)	,
(	34440	)	,
(	34425	)	,
(	34410	)	,
(	34395	)	,
(	34380	)	,
(	34365	)	,
(	34350	)	,
(	34335	)	,
(	34320	)	,
(	34305	)	,
(	34290	)	,
(	34275	)	,
(	34260	)	,
(	34245	)	,
(	34230	)	,
(	34215	)	,
(	34200	)	,
(	34185	)	,
(	34170	)	,
(	34155	)	,
(	34140	)	,
(	34125	)	,
(	34110	)	,
(	34095	)	,
(	34080	)	,
(	34065	)	,
(	34050	)	,
(	34035	)	,
(	34020	)	,
(	34005	)	,
(	33990	)	,
(	33975	)	,
(	33960	)	,
(	33945	)	,
(	33930	)	,
(	33915	)	,
(	33900	)	,
(	33885	)	,
(	33870	)	,
(	33855	)	,
(	33840	)	,
(	33825	)	,
(	33810	)	,
(	33795	)	,
(	33780	)	,
(	33765	)	,
(	33750	)	,
(	33735	)	,
(	33720	)	,
(	33705	)	,
(	33690	)	,
(	33675	)	,
(	33660	)	,
(	33645	)	,
(	33630	)	,
(	33615	)	,
(	33600	)	,
(	33585	)	,
(	33570	)	,
(	33555	)	,
(	33540	)	,
(	33525	)	,
(	33510	)	,
(	33495	)	,
(	33480	)	,
(	33465	)	,
(	33450	)	,
(	33435	)	,
(	33420	)	,
(	33405	)	,
(	33390	)	,
(	33375	)	,
(	33360	)	,
(	33345	)	,
(	33330	)	,
(	33315	)	,
(	33300	)	,
(	33285	)	,
(	33270	)	,
(	33255	)	,
(	33240	)	,
(	33225	)	,
(	33210	)	,
(	33195	)	,
(	33180	)	,
(	33165	)	,
(	33150	)	,
(	33135	)	,
(	33120	)	,
(	33105	)	,
(	33090	)	,
(	33075	)	,
(	33060	)	,
(	33045	)	,
(	33030	)	,
(	33015	)	,
(	33000	)	,
(	32985	)	,
(	32970	)	,
(	32955	)	,
(	32940	)	,
(	32925	)	,
(	32910	)	,
(	32895	)	,
(	32880	)	,
(	32865	)	,
(	32850	)	,
(	32835	)	,
(	32820	)	,
(	32805	)	,
(	32790	)	,
(	32775	)	,
(	32760	)	,
(	32745	)	,
(	32730	)	,
(	32715	)	,
(	32700	)	,
(	32685	)	,
(	32670	)	,
(	32655	)	,
(	32640	)	,
(	32625	)	,
(	32610	)	,
(	32595	)	,
(	32580	)	,
(	32565	)	,
(	32550	)	,
(	32535	)	,
(	32520	)	,
(	32505	)	,
(	32490	)	,
(	32475	)	,
(	32460	)	,
(	32445	)	,
(	32430	)	,
(	32415	)	,
(	32400	)	,
(	32385	)	,
(	32370	)	,
(	32355	)	,
(	32340	)	,
(	32325	)	,
(	32310	)	,
(	32295	)	,
(	32280	)	,
(	32265	)	,
(	32250	)	,
(	32235	)	,
(	32220	)	,
(	32205	)	,
(	32190	)	,
(	32175	)	,
(	32160	)	,
(	32145	)	,
(	32130	)	,
(	32115	)	,
(	32100	)	,
(	32085	)	,
(	32070	)	,
(	32055	)	,
(	32040	)	,
(	32025	)	,
(	32010	)	,
(	31995	)	,
(	31980	)	,
(	31965	)	,
(	31950	)	,
(	31935	)	,
(	31920	)	,
(	31905	)	,
(	31890	)	,
(	31875	)	,
(	31860	)	,
(	31845	)	,
(	31830	)	,
(	31815	)	,
(	31800	)	,
(	31785	)	,
(	31770	)	,
(	31755	)	,
(	31740	)	,
(	31725	)	,
(	31710	)	,
(	31695	)	,
(	31680	)	,
(	31665	)	,
(	31650	)	,
(	31635	)	,
(	31620	)	,
(	31605	)	,
(	31590	)	,
(	31575	)	,
(	31560	)	,
(	31545	)	,
(	31530	)	,
(	31515	)	,
(	31500	)	,
(	31485	)	,
(	31470	)	,
(	31455	)	,
(	31440	)	,
(	31425	)	,
(	31410	)	,
(	31395	)	,
(	31380	)	,
(	31365	)	,
(	31350	)	,
(	31335	)	,
(	31320	)	,
(	31305	)	,
(	31290	)	,
(	31275	)	,
(	31260	)	,
(	31245	)	,
(	31230	)	,
(	31215	)	,
(	31200	)	,
(	31185	)	,
(	31170	)	,
(	31155	)	,
(	31140	)	,
(	31125	)	,
(	31110	)	,
(	31095	)	,
(	31080	)	,
(	31065	)	,
(	31050	)	,
(	31035	)	,
(	31020	)	,
(	31005	)	,
(	30990	)	,
(	30975	)	,
(	30960	)	,
(	30945	)	,
(	30930	)	,
(	30915	)	,
(	30900	)	,
(	30885	)	,
(	30870	)	,
(	30855	)	,
(	30840	)	,
(	30825	)	,
(	30810	)	,
(	30795	)	,
(	30780	)	,
(	30765	)	,
(	30750	)	,
(	30735	)	,
(	30720	)	,
(	30705	)	,
(	30690	)	,
(	30675	)	,
(	30660	)	,
(	30645	)	,
(	30630	)	,
(	30615	)	,
(	30600	)	,
(	30585	)	,
(	30570	)	,
(	30555	)	,
(	30540	)	,
(	30525	)	,
(	30510	)	,
(	30495	)	,
(	30480	)	,
(	30465	)	,
(	30450	)	,
(	30435	)	,
(	30420	)	,
(	30405	)	,
(	30390	)	,
(	30375	)	,
(	30360	)	,
(	30345	)	,
(	30330	)	,
(	30315	)	,
(	30300	)	,
(	30285	)	,
(	30270	)	,
(	30255	)	,
(	30240	)	,
(	30225	)	,
(	30210	)	,
(	30195	)	,
(	30180	)	,
(	30165	)	,
(	30150	)	,
(	30135	)	,
(	30120	)	,
(	30105	)	,
(	30090	)	,
(	30075	)	,
(	30060	)	,
(	30045	)	,
(	30030	)	,
(	30015	)	,
(	30000	)	
 );
 
 end package LED_Flash_LUT_pkg;